--------------------------------------------------------------------------------
--                           IntAdder_16_f400_uid2
--                      (IntAdderClassical_16_f400_uid4)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_16_f400_uid2 is
   port ( XY : in  std_logic_vector(31 downto 0);
          --Y : in  std_logic_vector(15 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(31 downto 0)   );
end entity;

architecture arch of IntAdder_16_f400_uid2 is
begin
   --Classical
	R <= "0000000000000000" & ( XY(31 downto 16) + XY(15 downto 0) + Cin );
end architecture;

