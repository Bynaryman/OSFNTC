--------------------------------------------------------------------------------
--                  LZOCShifter_2_to_2_counting_4_F200_uid18
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: I OZb
-- Output signals: Count O

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZOCShifter_2_to_2_counting_4_F200_uid18 is
    port (clk : in std_logic;
          I : in  std_logic_vector(1 downto 0);
          OZb : in  std_logic;
          Count : out  std_logic_vector(1 downto 0);
          O : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of LZOCShifter_2_to_2_counting_4_F200_uid18 is
signal level2 :  std_logic_vector(1 downto 0);
signal sozb :  std_logic;
signal count1 :  std_logic;
signal level1 :  std_logic_vector(1 downto 0);
signal count0 :  std_logic;
signal level0 :  std_logic_vector(1 downto 0);
signal sCount :  std_logic_vector(1 downto 0);
begin
   level2 <= I ;
   sozb<= OZb;
   count1<= '1' when level2(1 downto 0) = (1 downto 0=>sozb) else '0';
   level1<= level2(1 downto 0) when count1='0' else (1 downto 0 => '0');

   count0<= '1' when level1(1 downto 1) = (1 downto 1=>sozb) else '0';
   level0<= level1(1 downto 0) when count0='0' else level1(0 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                                Arith_to_S3
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: BSC / UPC - Ledoux Louis
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: arith_i
-- Output signals: S3_o

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Arith_to_S3 is
    port (clk : in std_logic;
          arith_i : in  std_logic_vector(3 downto 0);
          S3_o : out  std_logic_vector(6 downto 0)   );
end entity;

architecture arch of Arith_to_S3 is
   component LZOCShifter_2_to_2_counting_4_F200_uid18 is
      port ( clk : in std_logic;
             I : in  std_logic_vector(1 downto 0);
             OZb : in  std_logic;
             Count : out  std_logic_vector(1 downto 0);
             O : out  std_logic_vector(1 downto 0)   );
   end component;

signal sign :  std_logic;
signal regime_check :  std_logic;
signal remainder :  std_logic_vector(1 downto 0);
signal not_s :  std_logic;
signal zero_NAR :  std_logic;
signal is_NAR :  std_logic;
signal implicit :  std_logic;
signal neg_count :  std_logic;
signal lzCount :  std_logic_vector(1 downto 0);
signal usefulBits :  std_logic_vector(1 downto 0);
signal extended_neg_count :  std_logic_vector(2 downto 0);
signal comp2_range_count :  std_logic_vector(2 downto 0);
signal fraction :  std_logic_vector(0 downto 0);
signal exponent :  std_logic_vector(2 downto 0);
signal biased_exponent :  std_logic_vector(2 downto 0);
begin
sign <= arith_i(3);
regime_check <= arith_i(2);
remainder <= arith_i(1 downto 0);
not_s <= not sign;
zero_NAR <= not regime_check when remainder="00" else '0';
is_NAR <= zero_NAR and sign;
implicit <= not(zero_NAR and not_s);
neg_count <= not (sign xor regime_check);
   lzoc: LZOCShifter_2_to_2_counting_4_F200_uid18
      port map ( clk  => clk,
                 I => remainder,
                 OZb => regime_check,
                 Count => lzCount,
                 O => usefulBits);
with neg_count  select  extended_neg_count <= 
   "111" when '1', 
   "000" when others;
comp2_range_count <= extended_neg_count xor ("0" & lzCount);
fraction <= usefulBits(0 downto 0);
exponent <= comp2_range_count;
biased_exponent <= exponent + 2;
S3_o <= is_NAR & sign & implicit & fraction & biased_exponent;
end architecture;

--------------------------------------------------------------------------------
--              LZOCShifterSticky_14_to_3_counting_16_F200_uid22
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: I OZb
-- Output signals: Count O Sticky

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZOCShifterSticky_14_to_3_counting_16_F200_uid22 is
    port (clk : in std_logic;
          I : in  std_logic_vector(13 downto 0);
          OZb : in  std_logic;
          Count : out  std_logic_vector(3 downto 0);
          O : out  std_logic_vector(2 downto 0);
          Sticky : out  std_logic   );
end entity;

architecture arch of LZOCShifterSticky_14_to_3_counting_16_F200_uid22 is
signal level4 :  std_logic_vector(13 downto 0);
signal sozb :  std_logic;
signal sticky4 :  std_logic;
signal count3 :  std_logic;
signal level3 :  std_logic_vector(13 downto 0);
signal sticky_high_3 :  std_logic;
signal sticky_low_3 :  std_logic;
signal sticky3 :  std_logic;
signal count2 :  std_logic;
signal level2 :  std_logic_vector(6 downto 0);
signal sticky_high_2 :  std_logic;
signal sticky_low_2 :  std_logic;
signal sticky2 :  std_logic;
signal count1 :  std_logic;
signal level1 :  std_logic_vector(3 downto 0);
signal sticky_high_1 :  std_logic;
signal sticky_low_1 :  std_logic;
signal sticky1 :  std_logic;
signal count0 :  std_logic;
signal level0 :  std_logic_vector(2 downto 0);
signal sticky_high_0 :  std_logic;
signal sticky_low_0 :  std_logic;
signal sticky0 :  std_logic;
signal sCount :  std_logic_vector(3 downto 0);
begin
   level4 <= I ;
   sozb<= OZb;
   sticky4 <= '0' ;
   count3<= '1' when level4(13 downto 6) = (13 downto 6=>sozb) else '0';
   level3<= level4(13 downto 0) when count3='0' else level4(5 downto 0) & (7 downto 0 => '0');
   sticky_high_3<= '0';
   sticky_low_3<= '0';
   sticky3<= sticky4 or sticky_high_3 when count3='0' else sticky4 or sticky_low_3;

   count2<= '1' when level3(13 downto 10) = (13 downto 10=>sozb) else '0';
   level2<= level3(13 downto 7) when count2='0' else level3(9 downto 3);
   sticky_high_2<= '0'when level3(6 downto 0) = CONV_STD_LOGIC_VECTOR(0,7) else '1';
   sticky_low_2<= '0'when level3(2 downto 0) = CONV_STD_LOGIC_VECTOR(0,3) else '1';
   sticky2<= sticky3 or sticky_high_2 when count2='0' else sticky3 or sticky_low_2;

   count1<= '1' when level2(6 downto 5) = (6 downto 5=>sozb) else '0';
   level1<= level2(6 downto 3) when count1='0' else level2(4 downto 1);
   sticky_high_1<= '0'when level2(2 downto 0) = CONV_STD_LOGIC_VECTOR(0,3) else '1';
   sticky_low_1<= '0'when level2(0 downto 0) = CONV_STD_LOGIC_VECTOR(0,1) else '1';
   sticky1<= sticky2 or sticky_high_1 when count1='0' else sticky2 or sticky_low_1;

   count0<= '1' when level1(3 downto 3) = (3 downto 3=>sozb) else '0';
   level0<= level1(3 downto 1) when count0='0' else level1(2 downto 0);
   sticky_high_0<= '0'when level1(0 downto 0) = CONV_STD_LOGIC_VECTOR(0,1) else '1';
   sticky_low_0<= '0';
   sticky0<= sticky1 or sticky_high_0 when count0='0' else sticky1 or sticky_low_0;

   O <= level0;
   sCount <= count3 & count2 & count1 & count0;
   Count <= sCount;
   Sticky <= sticky0;
end architecture;

--------------------------------------------------------------------------------
--                  RightShifterSticky4_by_max_4_F200_uid24
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X S padBit
-- Output signals: R Sticky

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity RightShifterSticky4_by_max_4_F200_uid24 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          S : in  std_logic_vector(2 downto 0);
          padBit : in  std_logic;
          R : out  std_logic_vector(3 downto 0);
          Sticky : out  std_logic   );
end entity;

architecture arch of RightShifterSticky4_by_max_4_F200_uid24 is
signal ps :  std_logic_vector(2 downto 0);
signal level3 :  std_logic_vector(3 downto 0);
signal stk2 :  std_logic;
signal level2 :  std_logic_vector(3 downto 0);
signal stk1 :  std_logic;
signal level1 :  std_logic_vector(3 downto 0);
signal stk0 :  std_logic;
signal level0 :  std_logic_vector(3 downto 0);
begin
   ps<= S;
   level3<= X;
   stk2 <= '1' when (level3(3 downto 0)/="0000" and ps(2)='1')   else '0';
   level2 <=  level3 when  ps(2)='0'    else (3 downto 0 => padBit) ;
   stk1 <= '1' when (level2(1 downto 0)/="00" and ps(1)='1') or stk2 ='1'   else '0';
   level1 <=  level2 when  ps(1)='0'    else (1 downto 0 => padBit) & level2(3 downto 2);
   stk0 <= '1' when (level1(0 downto 0)/="0" and ps(0)='1') or stk1 ='1'   else '0';
   level0 <=  level1 when  ps(0)='0'    else (0 downto 0 => padBit) & level1(3 downto 1);
   R <= level0;
   Sticky <= stk0;
end architecture;

--------------------------------------------------------------------------------
--                                    l2a
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Ledoux Louis - BSC / UPC
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: A isNaN
-- Output signals: arith_o

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity l2a is
    port (clk : in std_logic;
          A : in  std_logic_vector(13 downto 0);
          isNaN : in  std_logic;
          arith_o : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of l2a is
   component LZOCShifterSticky_14_to_3_counting_16_F200_uid22 is
      port ( clk : in std_logic;
             I : in  std_logic_vector(13 downto 0);
             OZb : in  std_logic;
             Count : out  std_logic_vector(3 downto 0);
             O : out  std_logic_vector(2 downto 0);
             Sticky : out  std_logic   );
   end component;

   component RightShifterSticky4_by_max_4_F200_uid24 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             S : in  std_logic_vector(2 downto 0);
             padBit : in  std_logic;
             R : out  std_logic_vector(3 downto 0);
             Sticky : out  std_logic   );
   end component;

signal rippled_carry :  std_logic_vector(13 downto 0);
signal count_bit, count_bit_d1 :  std_logic;
signal count_lzoc_o :  std_logic_vector(3 downto 0);
signal frac_lzoc_o :  std_logic_vector(2 downto 0);
signal sticky_lzoc_o :  std_logic;
signal unbiased_exp :  std_logic_vector(3 downto 0);
signal fraction :  std_logic_vector(1 downto 0);
signal bin_regime :  std_logic_vector(2 downto 0);
signal first_regime :  std_logic;
signal regime :  std_logic_vector(2 downto 0);
signal pad :  std_logic;
signal start_regime :  std_logic_vector(1 downto 0);
signal in_shift :  std_logic_vector(3 downto 0);
signal extended_posit :  std_logic_vector(3 downto 0);
signal pre_sticky :  std_logic;
signal truncated_posit, truncated_posit_d1 :  std_logic_vector(2 downto 0);
signal lsb :  std_logic;
signal guard :  std_logic;
signal sticky :  std_logic;
signal round_bit, round_bit_d1 :  std_logic;
signal is_NAR, is_NAR_d1 :  std_logic;
signal rounded_reg_exp_frac :  std_logic_vector(2 downto 0);
signal rounded_posit :  std_logic_vector(3 downto 0);
signal is_zero, is_zero_d1 :  std_logic;
signal rounded_posit_zero :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count_bit_d1 <=  count_bit;
            truncated_posit_d1 <=  truncated_posit;
            round_bit_d1 <=  round_bit;
            is_NAR_d1 <=  is_NAR;
            is_zero_d1 <=  is_zero;
         end if;
      end process;

   rippled_carry <= A;

--------------- Count 0/1 while shifting and sticky computation ---------------
   count_bit <= rippled_carry(13);
   lzoc_inst: LZOCShifterSticky_14_to_3_counting_16_F200_uid22
      port map ( clk  => clk,
                 I => rippled_carry,
                 OZb => count_bit,
                 Count => count_lzoc_o,
                 O => frac_lzoc_o,
                 Sticky => sticky_lzoc_o);

----------- Compute unbiased exponent from msb weigth and lzoc count -----------
   unbiased_exp <= CONV_STD_LOGIC_VECTOR(9,4) - (count_lzoc_o);
   fraction <= frac_lzoc_o (1 downto 0);
bin_regime<= unbiased_exp(2 downto 0);
first_regime<= unbiased_exp(3);
with first_regime  select  regime <= 
   bin_regime when '0', 
   not bin_regime when others;
pad<= not(first_regime xor count_bit);
with pad  select  start_regime <= 
   "01" when '0', 
   "10" when others; 
in_shift <= start_regime & fraction;
   rshift: RightShifterSticky4_by_max_4_F200_uid24
      port map ( clk  => clk,
                 S => regime,
                 X => in_shift,
                 padBit => pad,
                 R => extended_posit,
                 Sticky => pre_sticky);
truncated_posit<= extended_posit(3 downto 1);
lsb <= extended_posit(1);
guard <= extended_posit(0);
sticky <= fraction(0) or pre_sticky or sticky_lzoc_o;
round_bit<= guard and (sticky or lsb);
is_NAR<= isNaN;
rounded_reg_exp_frac<= truncated_posit_d1 + round_bit_d1;
rounded_posit <= count_bit_d1 & rounded_reg_exp_frac;
is_zero <= count_lzoc_o(3) when fraction="00" else '0';
rounded_posit_zero<= rounded_posit when is_zero_d1= '0' else "0000";
arith_o <= rounded_posit_zero when is_NAR_d1 = '0' else "1000";
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_2x2_F200_uid35
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_2x2_F200_uid35 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of DSPBlock_2x2_F200_uid35 is
signal Mint :  std_logic_vector(3 downto 0);
signal M :  std_logic_vector(3 downto 0);
signal Rtmp :  std_logic_vector(3 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(3 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          IntMultiplier_F200_uid31
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_F200_uid31 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplier_F200_uid31 is
   component DSPBlock_2x2_F200_uid35 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

signal XX_m32 :  std_logic_vector(1 downto 0);
signal YY_m32 :  std_logic_vector(1 downto 0);
signal tile_0_X :  std_logic_vector(1 downto 0);
signal tile_0_Y :  std_logic_vector(1 downto 0);
signal tile_0_output :  std_logic_vector(3 downto 0);
signal tile_0_filtered_output :  std_logic_vector(3 downto 0);
signal bh33_w0_0 :  std_logic;
signal bh33_w1_0 :  std_logic;
signal bh33_w2_0 :  std_logic;
signal bh33_w3_0 :  std_logic;
signal tmp_bitheapResult_bh33_3 :  std_logic_vector(3 downto 0);
signal bitheapResult_bh33 :  std_logic_vector(3 downto 0);
begin
   XX_m32 <= X ;
   YY_m32 <= Y ;
   tile_0_X <= X(1 downto 0);
   tile_0_Y <= Y(1 downto 0);
   tile_0_mult: DSPBlock_2x2_F200_uid35
      port map ( clk  => clk,
                 X => tile_0_X,
                 Y => tile_0_Y,
                 R => tile_0_output);

tile_0_filtered_output <= tile_0_output(3 downto 0);
   bh33_w0_0 <= tile_0_filtered_output(0);
   bh33_w1_0 <= tile_0_filtered_output(1);
   bh33_w2_0 <= tile_0_filtered_output(2);
   bh33_w3_0 <= tile_0_filtered_output(3);

   -- Adding the constant bits
      -- All the constant bits are zero, nothing to add

   tmp_bitheapResult_bh33_3 <= bh33_w3_0 & bh33_w2_0 & bh33_w1_0 & bh33_w0_0;
   bitheapResult_bh33 <= tmp_bitheapResult_bh33_3;
   R <= bitheapResult_bh33(3 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                     LeftShifter4_by_max_15_F200_uid38
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X S padBit
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter4_by_max_15_F200_uid38 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          S : in  std_logic_vector(3 downto 0);
          padBit : in  std_logic;
          R : out  std_logic_vector(18 downto 0)   );
end entity;

architecture arch of LeftShifter4_by_max_15_F200_uid38 is
signal ps :  std_logic_vector(3 downto 0);
signal level0 :  std_logic_vector(3 downto 0);
signal level1 :  std_logic_vector(4 downto 0);
signal level2 :  std_logic_vector(6 downto 0);
signal level3 :  std_logic_vector(10 downto 0);
signal level4 :  std_logic_vector(18 downto 0);
begin
   ps<= S;
   level0<= X;
   level1<= level0 & (0 downto 0 => '0') when ps(0)= '1' else     (0 downto 0 => padBit) & level0;
   level2<= level1 & (1 downto 0 => '0') when ps(1)= '1' else     (1 downto 0 => padBit) & level1;
   level3<= level2 & (3 downto 0 => '0') when ps(2)= '1' else     (3 downto 0 => padBit) & level2;
   level4<= level3 & (7 downto 0 => '0') when ps(3)= '1' else     (7 downto 0 => padBit) & level3;
   R <= level4(18 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                                   s3fdp
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Ledoux Louis - BSC / UPC
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: S3_x S3_y FTZ EOB
-- Output signals: A EOB_Q isNaN

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity s3fdp is
    port (clk, rst : in std_logic;
          S3_x : in  std_logic_vector(6 downto 0);
          S3_y : in  std_logic_vector(6 downto 0);
          FTZ : in  std_logic;
          EOB : in  std_logic;
          A : out  std_logic_vector(13 downto 0);
          EOB_Q : out  std_logic;
          isNaN : out  std_logic   );
end entity;

architecture arch of s3fdp is
   component IntMultiplier_F200_uid31 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component LeftShifter4_by_max_15_F200_uid38 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             S : in  std_logic_vector(3 downto 0);
             padBit : in  std_logic;
             R : out  std_logic_vector(18 downto 0)   );
   end component;

signal sign_X :  std_logic;
signal sign_Y :  std_logic;
signal sign_M :  std_logic;
signal isNaN_X :  std_logic;
signal isNaN_Y :  std_logic;
signal isNaN_M :  std_logic;
signal significand_X :  std_logic_vector(1 downto 0);
signal significand_Y :  std_logic_vector(1 downto 0);
signal significand_product :  std_logic_vector(3 downto 0);
signal scale_X_biased :  std_logic_vector(2 downto 0);
signal scale_Y_biased :  std_logic_vector(2 downto 0);
signal scale_product_twice_biased :  std_logic_vector(3 downto 0);
signal significand_product_cpt1 :  std_logic_vector(3 downto 0);
signal shift_value :  std_logic_vector(3 downto 0);
signal shifted_significand :  std_logic_vector(18 downto 0);
signal too_small :  std_logic;
signal too_big :  std_logic;
signal ext_summand1c :  std_logic_vector(13 downto 0);
signal not_ftz :  std_logic;
signal EOB_internal, EOB_internal_d1 :  std_logic;
signal not_ftz_sync :  std_logic;
signal carry_0_sync :  std_logic;
signal EOB_internal_delayed :  std_logic;
signal isNaN_M_sync :  std_logic;
signal too_big_sync :  std_logic;
signal isNaN_o, isNaN_o_d1 :  std_logic;
signal isNaN_delayed :  std_logic;
signal carry_0 :  std_logic;
signal summand_0 :  std_logic_vector(13 downto 0);
signal summand_and_carry_0 :  std_logic_vector(14 downto 0);
signal acc_0, acc_0_d1 :  std_logic_vector(14 downto 0);
signal acc_0_q :  std_logic_vector(14 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            EOB_internal_d1 <=  EOB_internal;
         end if;
      end process;
   process(clk, rst)
      begin
         if rst = '1' then
            isNaN_o_d1 <=  '0';
            acc_0_d1 <=  (others => '0');
         elsif clk'event and clk = '1' then
            isNaN_o_d1 <=  isNaN_o;
            acc_0_d1 <=  acc_0;
         end if;
      end process;
--------------------------- sign product processing ---------------------------
   sign_X <= S3_x(5);
   sign_Y <= S3_y(5);
   sign_M <= sign_X xor sign_Y;

---------------------------- NaN product processing ----------------------------
   isNaN_X <= S3_x(6);
   isNaN_Y <= S3_y(6);
   isNaN_M <= isNaN_X or isNaN_Y;

---------------------------- significand processing ----------------------------
   significand_X <= S3_x(4 downto 3);
   significand_Y <= S3_y(4 downto 3);
   significand_product_inst: IntMultiplier_F200_uid31
      port map ( clk  => clk,
                 X => significand_X,
                 Y => significand_Y,
                 R => significand_product);

------------------------------- scale processing -------------------------------
   scale_X_biased <= S3_x(2 downto 0);
   scale_Y_biased <= S3_y(2 downto 0);
   scale_product_twice_biased <= ("0" & scale_X_biased) + ("0" & scale_Y_biased);

--------------------------- pre-shift xoring (cpt1) ---------------------------
   significand_product_cpt1 <= significand_product when sign_M='0' else not(significand_product);

------------------------- significand product shifting -------------------------
   shift_value <= (scale_product_twice_biased) - (-1);
   significand_product_shifter_inst: LeftShifter4_by_max_15_F200_uid38
      port map ( clk  => clk,
                 S => shift_value,
                 X => significand_product_cpt1,
                 padBit => sign_M,
                 R => shifted_significand);

-------------- detect too low scale for this specific scratchpad --------------
   too_small <= '1' when (shift_value(3)='1') else '0';

-------------- detect too big scale for this specific scratchpad --------------
   too_big <= '1' when (unsigned(shift_value) > 8 and too_small='0') else '0';

--------------- shifted significand part select to form summand ---------------
   ext_summand1c <= "00000000000000" when too_small='1' else shifted_significand(16 downto 3);
----------------------------- Syncing some signals -----------------------------
   not_ftz <= not FTZ;
   EOB_internal <= EOB;
   not_ftz_sync <= not_ftz;
   carry_0_sync <= sign_M;
   EOB_internal_delayed <= EOB_internal_d1;
   isNaN_M_sync <= isNaN_M;
   too_big_sync <= too_big;

------------------------------ Output isNaN latch ------------------------------
   isNaN_o <= (too_big_sync or isNaN_M_sync or isNaN_delayed) when not_ftz_sync='1' else '0';
   isNaN_delayed <= isNaN_o_d1;

---------------------------- Carry Save Accumulator ----------------------------
   -- DQ logic
   acc_0_q <= acc_0_d1;

   -- sequential addition logic
   carry_0 <= carry_0_sync;
   summand_0 <= ext_summand1c(13 downto 0);
   summand_and_carry_0 <= ("0" & summand_0) + carry_0;
   acc_0 <= (("0" & acc_0_q(13 downto 0)) + summand_and_carry_0) when (not_ftz_sync='1') else
            summand_and_carry_0;

-------------------------------- Output Compose --------------------------------
   A <= acc_0_q(13 downto 0);

   EOB_Q <= EOB_internal_delayed;
   isNaN <= isNaN_delayed;
end architecture;

--------------------------------------------------------------------------------
--                                   PE_S3
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Ledoux Louis - BSC / UPC
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: s3_row_i_A s3_col_j_B C_out SOB EOB
-- Output signals: s3_row_im1_A s3_col_jm1_B SOB_Q EOB_Q C_out_Q

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity PE_S3 is
    port (clk, rst : in std_logic;
          s3_row_i_A : in  std_logic_vector(6 downto 0);
          s3_col_j_B : in  std_logic_vector(6 downto 0);
          C_out : in  std_logic_vector(14 downto 0);
          SOB : in  std_logic;
          EOB : in  std_logic;
          s3_row_im1_A : out  std_logic_vector(6 downto 0);
          s3_col_jm1_B : out  std_logic_vector(6 downto 0);
          SOB_Q : out  std_logic;
          EOB_Q : out  std_logic;
          C_out_Q : out  std_logic_vector(14 downto 0)   );
end entity;

architecture arch of PE_S3 is
   component s3fdp is
      port ( clk, rst : in std_logic;
             S3_x : in  std_logic_vector(6 downto 0);
             S3_y : in  std_logic_vector(6 downto 0);
             FTZ : in  std_logic;
             EOB : in  std_logic;
             A : out  std_logic_vector(13 downto 0);
             EOB_Q : out  std_logic;
             isNaN : out  std_logic   );
   end component;

signal s3_row_i_A_q :  std_logic_vector(6 downto 0);
signal s3_col_j_B_q :  std_logic_vector(6 downto 0);
signal sob_delayed :  std_logic;
signal eob_delayed :  std_logic;
signal mux_C_out, mux_C_out_d1, mux_C_out_d2 :  std_logic_vector(14 downto 0);
signal mux_C_out_HSSD :  std_logic_vector(14 downto 0);
signal isNaN_s3fdp :  std_logic;
signal EOB_s3fdp :  std_logic;
signal A_s3fdp :  std_logic_vector(13 downto 0);
signal s3_row_i_A_d1 :  std_logic_vector(6 downto 0);
signal s3_col_j_B_d1 :  std_logic_vector(6 downto 0);
signal SOB_d1 :  std_logic;
signal EOB_d1 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            mux_C_out_d1 <=  mux_C_out;
            mux_C_out_d2 <=  mux_C_out_d1;
            s3_row_i_A_d1 <=  s3_row_i_A;
            s3_col_j_B_d1 <=  s3_col_j_B;
            SOB_d1 <=  SOB;
            EOB_d1 <=  EOB;
         end if;
      end process;
------------------------ Functional delay z-1 of inputs ------------------------
   s3_row_i_A_q <= s3_row_i_A_d1;
   s3_col_j_B_q <= s3_col_j_B_d1;

------------------------- DQ flip flop for SOB and EOB -------------------------
   sob_delayed <= SOB_d1;
   eob_delayed <= EOB_d1;

----------------------------- Half Speed Sink Down -----------------------------
   with EOB_s3fdp  select  mux_C_out <= 
        (isNaN_s3fdp & A_s3fdp) when '1', 
        C_out when others;
   mux_C_out_HSSD <= mux_C_out_d2;

---------------------------- Instantiates the S3FDP ----------------------------
   s3fdp_inst: s3fdp
      port map ( clk => clk,
                 rst  => rst,
                 EOB => EOB,
                 FTZ => SOB,
                 S3_x => s3_row_i_A,
                 S3_y => s3_col_j_B,
                 A => A_s3fdp,
                 EOB_Q => EOB_s3fdp,
                 isNaN => isNaN_s3fdp);

------------------------- Compose the outputs signals -------------------------
   s3_row_im1_A <= s3_row_i_A_q;
   s3_col_jm1_B <= s3_col_j_B_q;
   SOB_Q <= sob_delayed;
   EOB_Q <= eob_delayed;
   C_out_Q <= mux_C_out_HSSD;
end architecture;

--------------------------------------------------------------------------------
--                            SystolicArrayKernel
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Ledoux Louis - BSC / UPC
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: rowsA colsB SOB EOB
-- Output signals: colsC EOB_Q_o

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity SystolicArrayKernel is
    port (clk, rst : in std_logic;
          rowsA : in  std_logic_vector(223 downto 0);
          colsB : in  std_logic_vector(216 downto 0);
          SOB : in  std_logic;
          EOB : in  std_logic;
          colsC : out  std_logic_vector(464 downto 0);
          EOB_Q_o : out  std_logic   );
end entity;

architecture arch of SystolicArrayKernel is
   component PE_S3 is
      port ( clk, rst : in std_logic;
             s3_row_i_A : in  std_logic_vector(6 downto 0);
             s3_col_j_B : in  std_logic_vector(6 downto 0);
             C_out : in  std_logic_vector(14 downto 0);
             SOB : in  std_logic;
             EOB : in  std_logic;
             s3_row_im1_A : out  std_logic_vector(6 downto 0);
             s3_col_jm1_B : out  std_logic_vector(6 downto 0);
             SOB_Q : out  std_logic;
             EOB_Q : out  std_logic;
             C_out_Q : out  std_logic_vector(14 downto 0)   );
   end component;

type T_2D_LAICPT2_np1_m is array(32 downto 0, 30 downto 0) of std_logic_vector(14 downto 0);
type T_2D_n_mp1 is array(31 downto 0, 31 downto 0) of std_logic_vector(6 downto 0);
type T_2D_np1_m is array(32 downto 0, 30 downto 0) of std_logic_vector(6 downto 0);
type T_2D_np1_m_logic is array(32 downto 0, 30 downto 0) of std_logic;
signal systolic_wires_rows_2D : T_2D_n_mp1;
signal systolic_wires_cols_2D : T_2D_np1_m;
signal systolic_sob_2D : T_2D_np1_m_logic;
signal systolic_eob_2D : T_2D_np1_m_logic;
signal systolic_C_out_2D : T_2D_LAICPT2_np1_m;
begin

----------------- Connect bus of B columns to top edges SA PEs -----------------
   cols_in: for JJ in 0 to 30 generate
      systolic_wires_cols_2D(0,JJ) <= colsB(((JJ+1)*7)-1 downto (JJ*7));
   end generate;

------------------ Connect bus of A rows to left edges SA PEs ------------------
   rows_in: for II in 0 to 31 generate
      systolic_wires_rows_2D(II,0) <= rowsA(((II+1)*7)-1 downto (II*7));
   end generate;

-------------- Connect the Start of Block signals of the TOP PEs --------------
   systolic_sob_2D(0,0) <= SOB;
   sob_1st_row: for JJ in 1 to 30 generate
      systolic_sob_2D(0,JJ) <= systolic_sob_2D(1,JJ-1);
   end generate;

--------------- Connect the End of Block signals of the TOP PEs ---------------
   systolic_eob_2D(0,0) <= EOB;
   eob_1st_row: for JJ in 1 to 30 generate
      systolic_eob_2D(0,JJ) <= systolic_eob_2D(1,JJ-1);
   end generate;

----------- Connect with 0s the input C carry out scheme of TOP PEs -----------
   C_out_input_1st_row: for JJ in 0 to 30 generate
      systolic_C_out_2D(0,JJ) <= "000000000000000";
   end generate;

------------------------- Connect PEs locally together -------------------------
   rows: for II in 0 to 31 generate
      cols: for JJ in 0 to 30 generate
         PE_ij: PE_S3
            port map ( clk => clk,
                       rst => rst,
                       s3_row_i_A => systolic_wires_rows_2D(II,JJ),
                       s3_col_j_B => systolic_wires_cols_2D(II,JJ),
                       SOB => systolic_sob_2D(II,JJ),
                       SOB_Q => systolic_sob_2D(II+1,JJ),
                       EOB => systolic_eob_2D(II,JJ),
                       EOB_Q => systolic_eob_2D(II+1,JJ),
                       C_out => systolic_C_out_2D(II,JJ),
                       C_out_Q => systolic_C_out_2D(II+1,JJ),
                       s3_row_im1_A => systolic_wires_rows_2D(II,JJ+1),
                       s3_col_jm1_B => systolic_wires_cols_2D(II+1,JJ));
      end generate;
   end generate;

------------------ Connect last row output C to output C bus ------------------
   cols_C_out: for JJ in 0 to 30 generate
      colsC(((JJ+1)*15)-1 downto (JJ*15)) <= systolic_C_out_2D(32,JJ);
   end generate;

------ Connect PE(N-1,M-1) EOB_Q to out world for valid data computation ------
   EOB_Q_o <= systolic_eob_2D(32,30);

end architecture;

--------------------------------------------------------------------------------
--                               SystolicArray
--              (SA_orthogonal_32w31h_posit_4_0_HSSD_F200_uid2)
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Ledoux Louis - BSC / UPC
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: rowsA colsB SOB EOB
-- Output signals: colsC EOB_Q_o

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity SystolicArray is
    port (clk, rst : in std_logic;
          rowsA : in  std_logic_vector(127 downto 0);
          colsB : in  std_logic_vector(123 downto 0);
          SOB : in  std_logic;
          EOB : in  std_logic;
          colsC : out  std_logic_vector(123 downto 0);
          EOB_Q_o : out  std_logic   );
end entity;

architecture arch of SystolicArray is
   component Arith_to_S3 is
      port ( clk : in std_logic;
             arith_i : in  std_logic_vector(3 downto 0);
             S3_o : out  std_logic_vector(6 downto 0)   );
   end component;

   component l2a is
      port ( clk : in std_logic;
             A : in  std_logic_vector(13 downto 0);
             isNaN : in  std_logic;
             arith_o : out  std_logic_vector(3 downto 0)   );
   end component;

   component SystolicArrayKernel is
      port ( clk, rst : in std_logic;
             rowsA : in  std_logic_vector(223 downto 0);
             colsB : in  std_logic_vector(216 downto 0);
             SOB : in  std_logic;
             EOB : in  std_logic;
             colsC : out  std_logic_vector(464 downto 0);
             EOB_Q_o : out  std_logic   );
   end component;

type array_M_dense is array(30 downto 0) of std_logic_vector(3 downto 0);
type array_M_s3 is array(30 downto 0) of std_logic_vector(6 downto 0);
type array_N_dense is array(31 downto 0) of std_logic_vector(3 downto 0);
type array_N_s3 is array(31 downto 0) of std_logic_vector(6 downto 0);
signal arith_in_row_0 :  std_logic_vector(3 downto 0);
signal arith_in_row_0_q0 :  std_logic_vector(3 downto 0);
signal arith_in_row_1, arith_in_row_1_d1 :  std_logic_vector(3 downto 0);
signal arith_in_row_1_q1 :  std_logic_vector(3 downto 0);
signal arith_in_row_2, arith_in_row_2_d1, arith_in_row_2_d2 :  std_logic_vector(3 downto 0);
signal arith_in_row_2_q2 :  std_logic_vector(3 downto 0);
signal arith_in_row_3, arith_in_row_3_d1, arith_in_row_3_d2, arith_in_row_3_d3 :  std_logic_vector(3 downto 0);
signal arith_in_row_3_q3 :  std_logic_vector(3 downto 0);
signal arith_in_row_4, arith_in_row_4_d1, arith_in_row_4_d2, arith_in_row_4_d3, arith_in_row_4_d4 :  std_logic_vector(3 downto 0);
signal arith_in_row_4_q4 :  std_logic_vector(3 downto 0);
signal arith_in_row_5, arith_in_row_5_d1, arith_in_row_5_d2, arith_in_row_5_d3, arith_in_row_5_d4, arith_in_row_5_d5 :  std_logic_vector(3 downto 0);
signal arith_in_row_5_q5 :  std_logic_vector(3 downto 0);
signal arith_in_row_6, arith_in_row_6_d1, arith_in_row_6_d2, arith_in_row_6_d3, arith_in_row_6_d4, arith_in_row_6_d5, arith_in_row_6_d6 :  std_logic_vector(3 downto 0);
signal arith_in_row_6_q6 :  std_logic_vector(3 downto 0);
signal arith_in_row_7, arith_in_row_7_d1, arith_in_row_7_d2, arith_in_row_7_d3, arith_in_row_7_d4, arith_in_row_7_d5, arith_in_row_7_d6, arith_in_row_7_d7 :  std_logic_vector(3 downto 0);
signal arith_in_row_7_q7 :  std_logic_vector(3 downto 0);
signal arith_in_row_8, arith_in_row_8_d1, arith_in_row_8_d2, arith_in_row_8_d3, arith_in_row_8_d4, arith_in_row_8_d5, arith_in_row_8_d6, arith_in_row_8_d7, arith_in_row_8_d8 :  std_logic_vector(3 downto 0);
signal arith_in_row_8_q8 :  std_logic_vector(3 downto 0);
signal arith_in_row_9, arith_in_row_9_d1, arith_in_row_9_d2, arith_in_row_9_d3, arith_in_row_9_d4, arith_in_row_9_d5, arith_in_row_9_d6, arith_in_row_9_d7, arith_in_row_9_d8, arith_in_row_9_d9 :  std_logic_vector(3 downto 0);
signal arith_in_row_9_q9 :  std_logic_vector(3 downto 0);
signal arith_in_row_10, arith_in_row_10_d1, arith_in_row_10_d2, arith_in_row_10_d3, arith_in_row_10_d4, arith_in_row_10_d5, arith_in_row_10_d6, arith_in_row_10_d7, arith_in_row_10_d8, arith_in_row_10_d9, arith_in_row_10_d10 :  std_logic_vector(3 downto 0);
signal arith_in_row_10_q10 :  std_logic_vector(3 downto 0);
signal arith_in_row_11, arith_in_row_11_d1, arith_in_row_11_d2, arith_in_row_11_d3, arith_in_row_11_d4, arith_in_row_11_d5, arith_in_row_11_d6, arith_in_row_11_d7, arith_in_row_11_d8, arith_in_row_11_d9, arith_in_row_11_d10, arith_in_row_11_d11 :  std_logic_vector(3 downto 0);
signal arith_in_row_11_q11 :  std_logic_vector(3 downto 0);
signal arith_in_row_12, arith_in_row_12_d1, arith_in_row_12_d2, arith_in_row_12_d3, arith_in_row_12_d4, arith_in_row_12_d5, arith_in_row_12_d6, arith_in_row_12_d7, arith_in_row_12_d8, arith_in_row_12_d9, arith_in_row_12_d10, arith_in_row_12_d11, arith_in_row_12_d12 :  std_logic_vector(3 downto 0);
signal arith_in_row_12_q12 :  std_logic_vector(3 downto 0);
signal arith_in_row_13, arith_in_row_13_d1, arith_in_row_13_d2, arith_in_row_13_d3, arith_in_row_13_d4, arith_in_row_13_d5, arith_in_row_13_d6, arith_in_row_13_d7, arith_in_row_13_d8, arith_in_row_13_d9, arith_in_row_13_d10, arith_in_row_13_d11, arith_in_row_13_d12, arith_in_row_13_d13 :  std_logic_vector(3 downto 0);
signal arith_in_row_13_q13 :  std_logic_vector(3 downto 0);
signal arith_in_row_14, arith_in_row_14_d1, arith_in_row_14_d2, arith_in_row_14_d3, arith_in_row_14_d4, arith_in_row_14_d5, arith_in_row_14_d6, arith_in_row_14_d7, arith_in_row_14_d8, arith_in_row_14_d9, arith_in_row_14_d10, arith_in_row_14_d11, arith_in_row_14_d12, arith_in_row_14_d13, arith_in_row_14_d14 :  std_logic_vector(3 downto 0);
signal arith_in_row_14_q14 :  std_logic_vector(3 downto 0);
signal arith_in_row_15, arith_in_row_15_d1, arith_in_row_15_d2, arith_in_row_15_d3, arith_in_row_15_d4, arith_in_row_15_d5, arith_in_row_15_d6, arith_in_row_15_d7, arith_in_row_15_d8, arith_in_row_15_d9, arith_in_row_15_d10, arith_in_row_15_d11, arith_in_row_15_d12, arith_in_row_15_d13, arith_in_row_15_d14, arith_in_row_15_d15 :  std_logic_vector(3 downto 0);
signal arith_in_row_15_q15 :  std_logic_vector(3 downto 0);
signal arith_in_row_16, arith_in_row_16_d1, arith_in_row_16_d2, arith_in_row_16_d3, arith_in_row_16_d4, arith_in_row_16_d5, arith_in_row_16_d6, arith_in_row_16_d7, arith_in_row_16_d8, arith_in_row_16_d9, arith_in_row_16_d10, arith_in_row_16_d11, arith_in_row_16_d12, arith_in_row_16_d13, arith_in_row_16_d14, arith_in_row_16_d15, arith_in_row_16_d16 :  std_logic_vector(3 downto 0);
signal arith_in_row_16_q16 :  std_logic_vector(3 downto 0);
signal arith_in_row_17, arith_in_row_17_d1, arith_in_row_17_d2, arith_in_row_17_d3, arith_in_row_17_d4, arith_in_row_17_d5, arith_in_row_17_d6, arith_in_row_17_d7, arith_in_row_17_d8, arith_in_row_17_d9, arith_in_row_17_d10, arith_in_row_17_d11, arith_in_row_17_d12, arith_in_row_17_d13, arith_in_row_17_d14, arith_in_row_17_d15, arith_in_row_17_d16, arith_in_row_17_d17 :  std_logic_vector(3 downto 0);
signal arith_in_row_17_q17 :  std_logic_vector(3 downto 0);
signal arith_in_row_18, arith_in_row_18_d1, arith_in_row_18_d2, arith_in_row_18_d3, arith_in_row_18_d4, arith_in_row_18_d5, arith_in_row_18_d6, arith_in_row_18_d7, arith_in_row_18_d8, arith_in_row_18_d9, arith_in_row_18_d10, arith_in_row_18_d11, arith_in_row_18_d12, arith_in_row_18_d13, arith_in_row_18_d14, arith_in_row_18_d15, arith_in_row_18_d16, arith_in_row_18_d17, arith_in_row_18_d18 :  std_logic_vector(3 downto 0);
signal arith_in_row_18_q18 :  std_logic_vector(3 downto 0);
signal arith_in_row_19, arith_in_row_19_d1, arith_in_row_19_d2, arith_in_row_19_d3, arith_in_row_19_d4, arith_in_row_19_d5, arith_in_row_19_d6, arith_in_row_19_d7, arith_in_row_19_d8, arith_in_row_19_d9, arith_in_row_19_d10, arith_in_row_19_d11, arith_in_row_19_d12, arith_in_row_19_d13, arith_in_row_19_d14, arith_in_row_19_d15, arith_in_row_19_d16, arith_in_row_19_d17, arith_in_row_19_d18, arith_in_row_19_d19 :  std_logic_vector(3 downto 0);
signal arith_in_row_19_q19 :  std_logic_vector(3 downto 0);
signal arith_in_row_20, arith_in_row_20_d1, arith_in_row_20_d2, arith_in_row_20_d3, arith_in_row_20_d4, arith_in_row_20_d5, arith_in_row_20_d6, arith_in_row_20_d7, arith_in_row_20_d8, arith_in_row_20_d9, arith_in_row_20_d10, arith_in_row_20_d11, arith_in_row_20_d12, arith_in_row_20_d13, arith_in_row_20_d14, arith_in_row_20_d15, arith_in_row_20_d16, arith_in_row_20_d17, arith_in_row_20_d18, arith_in_row_20_d19, arith_in_row_20_d20 :  std_logic_vector(3 downto 0);
signal arith_in_row_20_q20 :  std_logic_vector(3 downto 0);
signal arith_in_row_21, arith_in_row_21_d1, arith_in_row_21_d2, arith_in_row_21_d3, arith_in_row_21_d4, arith_in_row_21_d5, arith_in_row_21_d6, arith_in_row_21_d7, arith_in_row_21_d8, arith_in_row_21_d9, arith_in_row_21_d10, arith_in_row_21_d11, arith_in_row_21_d12, arith_in_row_21_d13, arith_in_row_21_d14, arith_in_row_21_d15, arith_in_row_21_d16, arith_in_row_21_d17, arith_in_row_21_d18, arith_in_row_21_d19, arith_in_row_21_d20, arith_in_row_21_d21 :  std_logic_vector(3 downto 0);
signal arith_in_row_21_q21 :  std_logic_vector(3 downto 0);
signal arith_in_row_22, arith_in_row_22_d1, arith_in_row_22_d2, arith_in_row_22_d3, arith_in_row_22_d4, arith_in_row_22_d5, arith_in_row_22_d6, arith_in_row_22_d7, arith_in_row_22_d8, arith_in_row_22_d9, arith_in_row_22_d10, arith_in_row_22_d11, arith_in_row_22_d12, arith_in_row_22_d13, arith_in_row_22_d14, arith_in_row_22_d15, arith_in_row_22_d16, arith_in_row_22_d17, arith_in_row_22_d18, arith_in_row_22_d19, arith_in_row_22_d20, arith_in_row_22_d21, arith_in_row_22_d22 :  std_logic_vector(3 downto 0);
signal arith_in_row_22_q22 :  std_logic_vector(3 downto 0);
signal arith_in_row_23, arith_in_row_23_d1, arith_in_row_23_d2, arith_in_row_23_d3, arith_in_row_23_d4, arith_in_row_23_d5, arith_in_row_23_d6, arith_in_row_23_d7, arith_in_row_23_d8, arith_in_row_23_d9, arith_in_row_23_d10, arith_in_row_23_d11, arith_in_row_23_d12, arith_in_row_23_d13, arith_in_row_23_d14, arith_in_row_23_d15, arith_in_row_23_d16, arith_in_row_23_d17, arith_in_row_23_d18, arith_in_row_23_d19, arith_in_row_23_d20, arith_in_row_23_d21, arith_in_row_23_d22, arith_in_row_23_d23 :  std_logic_vector(3 downto 0);
signal arith_in_row_23_q23 :  std_logic_vector(3 downto 0);
signal arith_in_row_24, arith_in_row_24_d1, arith_in_row_24_d2, arith_in_row_24_d3, arith_in_row_24_d4, arith_in_row_24_d5, arith_in_row_24_d6, arith_in_row_24_d7, arith_in_row_24_d8, arith_in_row_24_d9, arith_in_row_24_d10, arith_in_row_24_d11, arith_in_row_24_d12, arith_in_row_24_d13, arith_in_row_24_d14, arith_in_row_24_d15, arith_in_row_24_d16, arith_in_row_24_d17, arith_in_row_24_d18, arith_in_row_24_d19, arith_in_row_24_d20, arith_in_row_24_d21, arith_in_row_24_d22, arith_in_row_24_d23, arith_in_row_24_d24 :  std_logic_vector(3 downto 0);
signal arith_in_row_24_q24 :  std_logic_vector(3 downto 0);
signal arith_in_row_25, arith_in_row_25_d1, arith_in_row_25_d2, arith_in_row_25_d3, arith_in_row_25_d4, arith_in_row_25_d5, arith_in_row_25_d6, arith_in_row_25_d7, arith_in_row_25_d8, arith_in_row_25_d9, arith_in_row_25_d10, arith_in_row_25_d11, arith_in_row_25_d12, arith_in_row_25_d13, arith_in_row_25_d14, arith_in_row_25_d15, arith_in_row_25_d16, arith_in_row_25_d17, arith_in_row_25_d18, arith_in_row_25_d19, arith_in_row_25_d20, arith_in_row_25_d21, arith_in_row_25_d22, arith_in_row_25_d23, arith_in_row_25_d24, arith_in_row_25_d25 :  std_logic_vector(3 downto 0);
signal arith_in_row_25_q25 :  std_logic_vector(3 downto 0);
signal arith_in_row_26, arith_in_row_26_d1, arith_in_row_26_d2, arith_in_row_26_d3, arith_in_row_26_d4, arith_in_row_26_d5, arith_in_row_26_d6, arith_in_row_26_d7, arith_in_row_26_d8, arith_in_row_26_d9, arith_in_row_26_d10, arith_in_row_26_d11, arith_in_row_26_d12, arith_in_row_26_d13, arith_in_row_26_d14, arith_in_row_26_d15, arith_in_row_26_d16, arith_in_row_26_d17, arith_in_row_26_d18, arith_in_row_26_d19, arith_in_row_26_d20, arith_in_row_26_d21, arith_in_row_26_d22, arith_in_row_26_d23, arith_in_row_26_d24, arith_in_row_26_d25, arith_in_row_26_d26 :  std_logic_vector(3 downto 0);
signal arith_in_row_26_q26 :  std_logic_vector(3 downto 0);
signal arith_in_row_27, arith_in_row_27_d1, arith_in_row_27_d2, arith_in_row_27_d3, arith_in_row_27_d4, arith_in_row_27_d5, arith_in_row_27_d6, arith_in_row_27_d7, arith_in_row_27_d8, arith_in_row_27_d9, arith_in_row_27_d10, arith_in_row_27_d11, arith_in_row_27_d12, arith_in_row_27_d13, arith_in_row_27_d14, arith_in_row_27_d15, arith_in_row_27_d16, arith_in_row_27_d17, arith_in_row_27_d18, arith_in_row_27_d19, arith_in_row_27_d20, arith_in_row_27_d21, arith_in_row_27_d22, arith_in_row_27_d23, arith_in_row_27_d24, arith_in_row_27_d25, arith_in_row_27_d26, arith_in_row_27_d27 :  std_logic_vector(3 downto 0);
signal arith_in_row_27_q27 :  std_logic_vector(3 downto 0);
signal arith_in_row_28, arith_in_row_28_d1, arith_in_row_28_d2, arith_in_row_28_d3, arith_in_row_28_d4, arith_in_row_28_d5, arith_in_row_28_d6, arith_in_row_28_d7, arith_in_row_28_d8, arith_in_row_28_d9, arith_in_row_28_d10, arith_in_row_28_d11, arith_in_row_28_d12, arith_in_row_28_d13, arith_in_row_28_d14, arith_in_row_28_d15, arith_in_row_28_d16, arith_in_row_28_d17, arith_in_row_28_d18, arith_in_row_28_d19, arith_in_row_28_d20, arith_in_row_28_d21, arith_in_row_28_d22, arith_in_row_28_d23, arith_in_row_28_d24, arith_in_row_28_d25, arith_in_row_28_d26, arith_in_row_28_d27, arith_in_row_28_d28 :  std_logic_vector(3 downto 0);
signal arith_in_row_28_q28 :  std_logic_vector(3 downto 0);
signal arith_in_row_29, arith_in_row_29_d1, arith_in_row_29_d2, arith_in_row_29_d3, arith_in_row_29_d4, arith_in_row_29_d5, arith_in_row_29_d6, arith_in_row_29_d7, arith_in_row_29_d8, arith_in_row_29_d9, arith_in_row_29_d10, arith_in_row_29_d11, arith_in_row_29_d12, arith_in_row_29_d13, arith_in_row_29_d14, arith_in_row_29_d15, arith_in_row_29_d16, arith_in_row_29_d17, arith_in_row_29_d18, arith_in_row_29_d19, arith_in_row_29_d20, arith_in_row_29_d21, arith_in_row_29_d22, arith_in_row_29_d23, arith_in_row_29_d24, arith_in_row_29_d25, arith_in_row_29_d26, arith_in_row_29_d27, arith_in_row_29_d28, arith_in_row_29_d29 :  std_logic_vector(3 downto 0);
signal arith_in_row_29_q29 :  std_logic_vector(3 downto 0);
signal arith_in_row_30, arith_in_row_30_d1, arith_in_row_30_d2, arith_in_row_30_d3, arith_in_row_30_d4, arith_in_row_30_d5, arith_in_row_30_d6, arith_in_row_30_d7, arith_in_row_30_d8, arith_in_row_30_d9, arith_in_row_30_d10, arith_in_row_30_d11, arith_in_row_30_d12, arith_in_row_30_d13, arith_in_row_30_d14, arith_in_row_30_d15, arith_in_row_30_d16, arith_in_row_30_d17, arith_in_row_30_d18, arith_in_row_30_d19, arith_in_row_30_d20, arith_in_row_30_d21, arith_in_row_30_d22, arith_in_row_30_d23, arith_in_row_30_d24, arith_in_row_30_d25, arith_in_row_30_d26, arith_in_row_30_d27, arith_in_row_30_d28, arith_in_row_30_d29, arith_in_row_30_d30 :  std_logic_vector(3 downto 0);
signal arith_in_row_30_q30 :  std_logic_vector(3 downto 0);
signal arith_in_row_31, arith_in_row_31_d1, arith_in_row_31_d2, arith_in_row_31_d3, arith_in_row_31_d4, arith_in_row_31_d5, arith_in_row_31_d6, arith_in_row_31_d7, arith_in_row_31_d8, arith_in_row_31_d9, arith_in_row_31_d10, arith_in_row_31_d11, arith_in_row_31_d12, arith_in_row_31_d13, arith_in_row_31_d14, arith_in_row_31_d15, arith_in_row_31_d16, arith_in_row_31_d17, arith_in_row_31_d18, arith_in_row_31_d19, arith_in_row_31_d20, arith_in_row_31_d21, arith_in_row_31_d22, arith_in_row_31_d23, arith_in_row_31_d24, arith_in_row_31_d25, arith_in_row_31_d26, arith_in_row_31_d27, arith_in_row_31_d28, arith_in_row_31_d29, arith_in_row_31_d30, arith_in_row_31_d31 :  std_logic_vector(3 downto 0);
signal arith_in_row_31_q31 :  std_logic_vector(3 downto 0);
signal arith_in_col_0 :  std_logic_vector(3 downto 0);
signal arith_in_col_0_q0 :  std_logic_vector(3 downto 0);
signal arith_in_col_1, arith_in_col_1_d1 :  std_logic_vector(3 downto 0);
signal arith_in_col_1_q1 :  std_logic_vector(3 downto 0);
signal arith_in_col_2, arith_in_col_2_d1, arith_in_col_2_d2 :  std_logic_vector(3 downto 0);
signal arith_in_col_2_q2 :  std_logic_vector(3 downto 0);
signal arith_in_col_3, arith_in_col_3_d1, arith_in_col_3_d2, arith_in_col_3_d3 :  std_logic_vector(3 downto 0);
signal arith_in_col_3_q3 :  std_logic_vector(3 downto 0);
signal arith_in_col_4, arith_in_col_4_d1, arith_in_col_4_d2, arith_in_col_4_d3, arith_in_col_4_d4 :  std_logic_vector(3 downto 0);
signal arith_in_col_4_q4 :  std_logic_vector(3 downto 0);
signal arith_in_col_5, arith_in_col_5_d1, arith_in_col_5_d2, arith_in_col_5_d3, arith_in_col_5_d4, arith_in_col_5_d5 :  std_logic_vector(3 downto 0);
signal arith_in_col_5_q5 :  std_logic_vector(3 downto 0);
signal arith_in_col_6, arith_in_col_6_d1, arith_in_col_6_d2, arith_in_col_6_d3, arith_in_col_6_d4, arith_in_col_6_d5, arith_in_col_6_d6 :  std_logic_vector(3 downto 0);
signal arith_in_col_6_q6 :  std_logic_vector(3 downto 0);
signal arith_in_col_7, arith_in_col_7_d1, arith_in_col_7_d2, arith_in_col_7_d3, arith_in_col_7_d4, arith_in_col_7_d5, arith_in_col_7_d6, arith_in_col_7_d7 :  std_logic_vector(3 downto 0);
signal arith_in_col_7_q7 :  std_logic_vector(3 downto 0);
signal arith_in_col_8, arith_in_col_8_d1, arith_in_col_8_d2, arith_in_col_8_d3, arith_in_col_8_d4, arith_in_col_8_d5, arith_in_col_8_d6, arith_in_col_8_d7, arith_in_col_8_d8 :  std_logic_vector(3 downto 0);
signal arith_in_col_8_q8 :  std_logic_vector(3 downto 0);
signal arith_in_col_9, arith_in_col_9_d1, arith_in_col_9_d2, arith_in_col_9_d3, arith_in_col_9_d4, arith_in_col_9_d5, arith_in_col_9_d6, arith_in_col_9_d7, arith_in_col_9_d8, arith_in_col_9_d9 :  std_logic_vector(3 downto 0);
signal arith_in_col_9_q9 :  std_logic_vector(3 downto 0);
signal arith_in_col_10, arith_in_col_10_d1, arith_in_col_10_d2, arith_in_col_10_d3, arith_in_col_10_d4, arith_in_col_10_d5, arith_in_col_10_d6, arith_in_col_10_d7, arith_in_col_10_d8, arith_in_col_10_d9, arith_in_col_10_d10 :  std_logic_vector(3 downto 0);
signal arith_in_col_10_q10 :  std_logic_vector(3 downto 0);
signal arith_in_col_11, arith_in_col_11_d1, arith_in_col_11_d2, arith_in_col_11_d3, arith_in_col_11_d4, arith_in_col_11_d5, arith_in_col_11_d6, arith_in_col_11_d7, arith_in_col_11_d8, arith_in_col_11_d9, arith_in_col_11_d10, arith_in_col_11_d11 :  std_logic_vector(3 downto 0);
signal arith_in_col_11_q11 :  std_logic_vector(3 downto 0);
signal arith_in_col_12, arith_in_col_12_d1, arith_in_col_12_d2, arith_in_col_12_d3, arith_in_col_12_d4, arith_in_col_12_d5, arith_in_col_12_d6, arith_in_col_12_d7, arith_in_col_12_d8, arith_in_col_12_d9, arith_in_col_12_d10, arith_in_col_12_d11, arith_in_col_12_d12 :  std_logic_vector(3 downto 0);
signal arith_in_col_12_q12 :  std_logic_vector(3 downto 0);
signal arith_in_col_13, arith_in_col_13_d1, arith_in_col_13_d2, arith_in_col_13_d3, arith_in_col_13_d4, arith_in_col_13_d5, arith_in_col_13_d6, arith_in_col_13_d7, arith_in_col_13_d8, arith_in_col_13_d9, arith_in_col_13_d10, arith_in_col_13_d11, arith_in_col_13_d12, arith_in_col_13_d13 :  std_logic_vector(3 downto 0);
signal arith_in_col_13_q13 :  std_logic_vector(3 downto 0);
signal arith_in_col_14, arith_in_col_14_d1, arith_in_col_14_d2, arith_in_col_14_d3, arith_in_col_14_d4, arith_in_col_14_d5, arith_in_col_14_d6, arith_in_col_14_d7, arith_in_col_14_d8, arith_in_col_14_d9, arith_in_col_14_d10, arith_in_col_14_d11, arith_in_col_14_d12, arith_in_col_14_d13, arith_in_col_14_d14 :  std_logic_vector(3 downto 0);
signal arith_in_col_14_q14 :  std_logic_vector(3 downto 0);
signal arith_in_col_15, arith_in_col_15_d1, arith_in_col_15_d2, arith_in_col_15_d3, arith_in_col_15_d4, arith_in_col_15_d5, arith_in_col_15_d6, arith_in_col_15_d7, arith_in_col_15_d8, arith_in_col_15_d9, arith_in_col_15_d10, arith_in_col_15_d11, arith_in_col_15_d12, arith_in_col_15_d13, arith_in_col_15_d14, arith_in_col_15_d15 :  std_logic_vector(3 downto 0);
signal arith_in_col_15_q15 :  std_logic_vector(3 downto 0);
signal arith_in_col_16, arith_in_col_16_d1, arith_in_col_16_d2, arith_in_col_16_d3, arith_in_col_16_d4, arith_in_col_16_d5, arith_in_col_16_d6, arith_in_col_16_d7, arith_in_col_16_d8, arith_in_col_16_d9, arith_in_col_16_d10, arith_in_col_16_d11, arith_in_col_16_d12, arith_in_col_16_d13, arith_in_col_16_d14, arith_in_col_16_d15, arith_in_col_16_d16 :  std_logic_vector(3 downto 0);
signal arith_in_col_16_q16 :  std_logic_vector(3 downto 0);
signal arith_in_col_17, arith_in_col_17_d1, arith_in_col_17_d2, arith_in_col_17_d3, arith_in_col_17_d4, arith_in_col_17_d5, arith_in_col_17_d6, arith_in_col_17_d7, arith_in_col_17_d8, arith_in_col_17_d9, arith_in_col_17_d10, arith_in_col_17_d11, arith_in_col_17_d12, arith_in_col_17_d13, arith_in_col_17_d14, arith_in_col_17_d15, arith_in_col_17_d16, arith_in_col_17_d17 :  std_logic_vector(3 downto 0);
signal arith_in_col_17_q17 :  std_logic_vector(3 downto 0);
signal arith_in_col_18, arith_in_col_18_d1, arith_in_col_18_d2, arith_in_col_18_d3, arith_in_col_18_d4, arith_in_col_18_d5, arith_in_col_18_d6, arith_in_col_18_d7, arith_in_col_18_d8, arith_in_col_18_d9, arith_in_col_18_d10, arith_in_col_18_d11, arith_in_col_18_d12, arith_in_col_18_d13, arith_in_col_18_d14, arith_in_col_18_d15, arith_in_col_18_d16, arith_in_col_18_d17, arith_in_col_18_d18 :  std_logic_vector(3 downto 0);
signal arith_in_col_18_q18 :  std_logic_vector(3 downto 0);
signal arith_in_col_19, arith_in_col_19_d1, arith_in_col_19_d2, arith_in_col_19_d3, arith_in_col_19_d4, arith_in_col_19_d5, arith_in_col_19_d6, arith_in_col_19_d7, arith_in_col_19_d8, arith_in_col_19_d9, arith_in_col_19_d10, arith_in_col_19_d11, arith_in_col_19_d12, arith_in_col_19_d13, arith_in_col_19_d14, arith_in_col_19_d15, arith_in_col_19_d16, arith_in_col_19_d17, arith_in_col_19_d18, arith_in_col_19_d19 :  std_logic_vector(3 downto 0);
signal arith_in_col_19_q19 :  std_logic_vector(3 downto 0);
signal arith_in_col_20, arith_in_col_20_d1, arith_in_col_20_d2, arith_in_col_20_d3, arith_in_col_20_d4, arith_in_col_20_d5, arith_in_col_20_d6, arith_in_col_20_d7, arith_in_col_20_d8, arith_in_col_20_d9, arith_in_col_20_d10, arith_in_col_20_d11, arith_in_col_20_d12, arith_in_col_20_d13, arith_in_col_20_d14, arith_in_col_20_d15, arith_in_col_20_d16, arith_in_col_20_d17, arith_in_col_20_d18, arith_in_col_20_d19, arith_in_col_20_d20 :  std_logic_vector(3 downto 0);
signal arith_in_col_20_q20 :  std_logic_vector(3 downto 0);
signal arith_in_col_21, arith_in_col_21_d1, arith_in_col_21_d2, arith_in_col_21_d3, arith_in_col_21_d4, arith_in_col_21_d5, arith_in_col_21_d6, arith_in_col_21_d7, arith_in_col_21_d8, arith_in_col_21_d9, arith_in_col_21_d10, arith_in_col_21_d11, arith_in_col_21_d12, arith_in_col_21_d13, arith_in_col_21_d14, arith_in_col_21_d15, arith_in_col_21_d16, arith_in_col_21_d17, arith_in_col_21_d18, arith_in_col_21_d19, arith_in_col_21_d20, arith_in_col_21_d21 :  std_logic_vector(3 downto 0);
signal arith_in_col_21_q21 :  std_logic_vector(3 downto 0);
signal arith_in_col_22, arith_in_col_22_d1, arith_in_col_22_d2, arith_in_col_22_d3, arith_in_col_22_d4, arith_in_col_22_d5, arith_in_col_22_d6, arith_in_col_22_d7, arith_in_col_22_d8, arith_in_col_22_d9, arith_in_col_22_d10, arith_in_col_22_d11, arith_in_col_22_d12, arith_in_col_22_d13, arith_in_col_22_d14, arith_in_col_22_d15, arith_in_col_22_d16, arith_in_col_22_d17, arith_in_col_22_d18, arith_in_col_22_d19, arith_in_col_22_d20, arith_in_col_22_d21, arith_in_col_22_d22 :  std_logic_vector(3 downto 0);
signal arith_in_col_22_q22 :  std_logic_vector(3 downto 0);
signal arith_in_col_23, arith_in_col_23_d1, arith_in_col_23_d2, arith_in_col_23_d3, arith_in_col_23_d4, arith_in_col_23_d5, arith_in_col_23_d6, arith_in_col_23_d7, arith_in_col_23_d8, arith_in_col_23_d9, arith_in_col_23_d10, arith_in_col_23_d11, arith_in_col_23_d12, arith_in_col_23_d13, arith_in_col_23_d14, arith_in_col_23_d15, arith_in_col_23_d16, arith_in_col_23_d17, arith_in_col_23_d18, arith_in_col_23_d19, arith_in_col_23_d20, arith_in_col_23_d21, arith_in_col_23_d22, arith_in_col_23_d23 :  std_logic_vector(3 downto 0);
signal arith_in_col_23_q23 :  std_logic_vector(3 downto 0);
signal arith_in_col_24, arith_in_col_24_d1, arith_in_col_24_d2, arith_in_col_24_d3, arith_in_col_24_d4, arith_in_col_24_d5, arith_in_col_24_d6, arith_in_col_24_d7, arith_in_col_24_d8, arith_in_col_24_d9, arith_in_col_24_d10, arith_in_col_24_d11, arith_in_col_24_d12, arith_in_col_24_d13, arith_in_col_24_d14, arith_in_col_24_d15, arith_in_col_24_d16, arith_in_col_24_d17, arith_in_col_24_d18, arith_in_col_24_d19, arith_in_col_24_d20, arith_in_col_24_d21, arith_in_col_24_d22, arith_in_col_24_d23, arith_in_col_24_d24 :  std_logic_vector(3 downto 0);
signal arith_in_col_24_q24 :  std_logic_vector(3 downto 0);
signal arith_in_col_25, arith_in_col_25_d1, arith_in_col_25_d2, arith_in_col_25_d3, arith_in_col_25_d4, arith_in_col_25_d5, arith_in_col_25_d6, arith_in_col_25_d7, arith_in_col_25_d8, arith_in_col_25_d9, arith_in_col_25_d10, arith_in_col_25_d11, arith_in_col_25_d12, arith_in_col_25_d13, arith_in_col_25_d14, arith_in_col_25_d15, arith_in_col_25_d16, arith_in_col_25_d17, arith_in_col_25_d18, arith_in_col_25_d19, arith_in_col_25_d20, arith_in_col_25_d21, arith_in_col_25_d22, arith_in_col_25_d23, arith_in_col_25_d24, arith_in_col_25_d25 :  std_logic_vector(3 downto 0);
signal arith_in_col_25_q25 :  std_logic_vector(3 downto 0);
signal arith_in_col_26, arith_in_col_26_d1, arith_in_col_26_d2, arith_in_col_26_d3, arith_in_col_26_d4, arith_in_col_26_d5, arith_in_col_26_d6, arith_in_col_26_d7, arith_in_col_26_d8, arith_in_col_26_d9, arith_in_col_26_d10, arith_in_col_26_d11, arith_in_col_26_d12, arith_in_col_26_d13, arith_in_col_26_d14, arith_in_col_26_d15, arith_in_col_26_d16, arith_in_col_26_d17, arith_in_col_26_d18, arith_in_col_26_d19, arith_in_col_26_d20, arith_in_col_26_d21, arith_in_col_26_d22, arith_in_col_26_d23, arith_in_col_26_d24, arith_in_col_26_d25, arith_in_col_26_d26 :  std_logic_vector(3 downto 0);
signal arith_in_col_26_q26 :  std_logic_vector(3 downto 0);
signal arith_in_col_27, arith_in_col_27_d1, arith_in_col_27_d2, arith_in_col_27_d3, arith_in_col_27_d4, arith_in_col_27_d5, arith_in_col_27_d6, arith_in_col_27_d7, arith_in_col_27_d8, arith_in_col_27_d9, arith_in_col_27_d10, arith_in_col_27_d11, arith_in_col_27_d12, arith_in_col_27_d13, arith_in_col_27_d14, arith_in_col_27_d15, arith_in_col_27_d16, arith_in_col_27_d17, arith_in_col_27_d18, arith_in_col_27_d19, arith_in_col_27_d20, arith_in_col_27_d21, arith_in_col_27_d22, arith_in_col_27_d23, arith_in_col_27_d24, arith_in_col_27_d25, arith_in_col_27_d26, arith_in_col_27_d27 :  std_logic_vector(3 downto 0);
signal arith_in_col_27_q27 :  std_logic_vector(3 downto 0);
signal arith_in_col_28, arith_in_col_28_d1, arith_in_col_28_d2, arith_in_col_28_d3, arith_in_col_28_d4, arith_in_col_28_d5, arith_in_col_28_d6, arith_in_col_28_d7, arith_in_col_28_d8, arith_in_col_28_d9, arith_in_col_28_d10, arith_in_col_28_d11, arith_in_col_28_d12, arith_in_col_28_d13, arith_in_col_28_d14, arith_in_col_28_d15, arith_in_col_28_d16, arith_in_col_28_d17, arith_in_col_28_d18, arith_in_col_28_d19, arith_in_col_28_d20, arith_in_col_28_d21, arith_in_col_28_d22, arith_in_col_28_d23, arith_in_col_28_d24, arith_in_col_28_d25, arith_in_col_28_d26, arith_in_col_28_d27, arith_in_col_28_d28 :  std_logic_vector(3 downto 0);
signal arith_in_col_28_q28 :  std_logic_vector(3 downto 0);
signal arith_in_col_29, arith_in_col_29_d1, arith_in_col_29_d2, arith_in_col_29_d3, arith_in_col_29_d4, arith_in_col_29_d5, arith_in_col_29_d6, arith_in_col_29_d7, arith_in_col_29_d8, arith_in_col_29_d9, arith_in_col_29_d10, arith_in_col_29_d11, arith_in_col_29_d12, arith_in_col_29_d13, arith_in_col_29_d14, arith_in_col_29_d15, arith_in_col_29_d16, arith_in_col_29_d17, arith_in_col_29_d18, arith_in_col_29_d19, arith_in_col_29_d20, arith_in_col_29_d21, arith_in_col_29_d22, arith_in_col_29_d23, arith_in_col_29_d24, arith_in_col_29_d25, arith_in_col_29_d26, arith_in_col_29_d27, arith_in_col_29_d28, arith_in_col_29_d29 :  std_logic_vector(3 downto 0);
signal arith_in_col_29_q29 :  std_logic_vector(3 downto 0);
signal arith_in_col_30, arith_in_col_30_d1, arith_in_col_30_d2, arith_in_col_30_d3, arith_in_col_30_d4, arith_in_col_30_d5, arith_in_col_30_d6, arith_in_col_30_d7, arith_in_col_30_d8, arith_in_col_30_d9, arith_in_col_30_d10, arith_in_col_30_d11, arith_in_col_30_d12, arith_in_col_30_d13, arith_in_col_30_d14, arith_in_col_30_d15, arith_in_col_30_d16, arith_in_col_30_d17, arith_in_col_30_d18, arith_in_col_30_d19, arith_in_col_30_d20, arith_in_col_30_d21, arith_in_col_30_d22, arith_in_col_30_d23, arith_in_col_30_d24, arith_in_col_30_d25, arith_in_col_30_d26, arith_in_col_30_d27, arith_in_col_30_d28, arith_in_col_30_d29, arith_in_col_30_d30 :  std_logic_vector(3 downto 0);
signal arith_in_col_30_q30 :  std_logic_vector(3 downto 0);
signal colsC_LAICPT2 :  std_logic_vector(464 downto 0);
signal SOB_select :  std_logic;
signal SOB_q0 :  std_logic;
signal EOB_select :  std_logic;
signal EOB_q0 :  std_logic;
signal LAICPT2_to_arith :  std_logic_vector(123 downto 0);
signal arith_out_col_out_0, arith_out_col_out_0_d1, arith_out_col_out_0_d2, arith_out_col_out_0_d3, arith_out_col_out_0_d4, arith_out_col_out_0_d5, arith_out_col_out_0_d6, arith_out_col_out_0_d7, arith_out_col_out_0_d8, arith_out_col_out_0_d9, arith_out_col_out_0_d10, arith_out_col_out_0_d11, arith_out_col_out_0_d12, arith_out_col_out_0_d13, arith_out_col_out_0_d14, arith_out_col_out_0_d15, arith_out_col_out_0_d16, arith_out_col_out_0_d17, arith_out_col_out_0_d18, arith_out_col_out_0_d19, arith_out_col_out_0_d20, arith_out_col_out_0_d21, arith_out_col_out_0_d22, arith_out_col_out_0_d23, arith_out_col_out_0_d24, arith_out_col_out_0_d25, arith_out_col_out_0_d26, arith_out_col_out_0_d27, arith_out_col_out_0_d28, arith_out_col_out_0_d29, arith_out_col_out_0_d30 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_0_q30 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_1, arith_out_col_out_1_d1, arith_out_col_out_1_d2, arith_out_col_out_1_d3, arith_out_col_out_1_d4, arith_out_col_out_1_d5, arith_out_col_out_1_d6, arith_out_col_out_1_d7, arith_out_col_out_1_d8, arith_out_col_out_1_d9, arith_out_col_out_1_d10, arith_out_col_out_1_d11, arith_out_col_out_1_d12, arith_out_col_out_1_d13, arith_out_col_out_1_d14, arith_out_col_out_1_d15, arith_out_col_out_1_d16, arith_out_col_out_1_d17, arith_out_col_out_1_d18, arith_out_col_out_1_d19, arith_out_col_out_1_d20, arith_out_col_out_1_d21, arith_out_col_out_1_d22, arith_out_col_out_1_d23, arith_out_col_out_1_d24, arith_out_col_out_1_d25, arith_out_col_out_1_d26, arith_out_col_out_1_d27, arith_out_col_out_1_d28, arith_out_col_out_1_d29 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_1_q29 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_2, arith_out_col_out_2_d1, arith_out_col_out_2_d2, arith_out_col_out_2_d3, arith_out_col_out_2_d4, arith_out_col_out_2_d5, arith_out_col_out_2_d6, arith_out_col_out_2_d7, arith_out_col_out_2_d8, arith_out_col_out_2_d9, arith_out_col_out_2_d10, arith_out_col_out_2_d11, arith_out_col_out_2_d12, arith_out_col_out_2_d13, arith_out_col_out_2_d14, arith_out_col_out_2_d15, arith_out_col_out_2_d16, arith_out_col_out_2_d17, arith_out_col_out_2_d18, arith_out_col_out_2_d19, arith_out_col_out_2_d20, arith_out_col_out_2_d21, arith_out_col_out_2_d22, arith_out_col_out_2_d23, arith_out_col_out_2_d24, arith_out_col_out_2_d25, arith_out_col_out_2_d26, arith_out_col_out_2_d27, arith_out_col_out_2_d28 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_2_q28 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_3, arith_out_col_out_3_d1, arith_out_col_out_3_d2, arith_out_col_out_3_d3, arith_out_col_out_3_d4, arith_out_col_out_3_d5, arith_out_col_out_3_d6, arith_out_col_out_3_d7, arith_out_col_out_3_d8, arith_out_col_out_3_d9, arith_out_col_out_3_d10, arith_out_col_out_3_d11, arith_out_col_out_3_d12, arith_out_col_out_3_d13, arith_out_col_out_3_d14, arith_out_col_out_3_d15, arith_out_col_out_3_d16, arith_out_col_out_3_d17, arith_out_col_out_3_d18, arith_out_col_out_3_d19, arith_out_col_out_3_d20, arith_out_col_out_3_d21, arith_out_col_out_3_d22, arith_out_col_out_3_d23, arith_out_col_out_3_d24, arith_out_col_out_3_d25, arith_out_col_out_3_d26, arith_out_col_out_3_d27 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_3_q27 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_4, arith_out_col_out_4_d1, arith_out_col_out_4_d2, arith_out_col_out_4_d3, arith_out_col_out_4_d4, arith_out_col_out_4_d5, arith_out_col_out_4_d6, arith_out_col_out_4_d7, arith_out_col_out_4_d8, arith_out_col_out_4_d9, arith_out_col_out_4_d10, arith_out_col_out_4_d11, arith_out_col_out_4_d12, arith_out_col_out_4_d13, arith_out_col_out_4_d14, arith_out_col_out_4_d15, arith_out_col_out_4_d16, arith_out_col_out_4_d17, arith_out_col_out_4_d18, arith_out_col_out_4_d19, arith_out_col_out_4_d20, arith_out_col_out_4_d21, arith_out_col_out_4_d22, arith_out_col_out_4_d23, arith_out_col_out_4_d24, arith_out_col_out_4_d25, arith_out_col_out_4_d26 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_4_q26 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_5, arith_out_col_out_5_d1, arith_out_col_out_5_d2, arith_out_col_out_5_d3, arith_out_col_out_5_d4, arith_out_col_out_5_d5, arith_out_col_out_5_d6, arith_out_col_out_5_d7, arith_out_col_out_5_d8, arith_out_col_out_5_d9, arith_out_col_out_5_d10, arith_out_col_out_5_d11, arith_out_col_out_5_d12, arith_out_col_out_5_d13, arith_out_col_out_5_d14, arith_out_col_out_5_d15, arith_out_col_out_5_d16, arith_out_col_out_5_d17, arith_out_col_out_5_d18, arith_out_col_out_5_d19, arith_out_col_out_5_d20, arith_out_col_out_5_d21, arith_out_col_out_5_d22, arith_out_col_out_5_d23, arith_out_col_out_5_d24, arith_out_col_out_5_d25 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_5_q25 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_6, arith_out_col_out_6_d1, arith_out_col_out_6_d2, arith_out_col_out_6_d3, arith_out_col_out_6_d4, arith_out_col_out_6_d5, arith_out_col_out_6_d6, arith_out_col_out_6_d7, arith_out_col_out_6_d8, arith_out_col_out_6_d9, arith_out_col_out_6_d10, arith_out_col_out_6_d11, arith_out_col_out_6_d12, arith_out_col_out_6_d13, arith_out_col_out_6_d14, arith_out_col_out_6_d15, arith_out_col_out_6_d16, arith_out_col_out_6_d17, arith_out_col_out_6_d18, arith_out_col_out_6_d19, arith_out_col_out_6_d20, arith_out_col_out_6_d21, arith_out_col_out_6_d22, arith_out_col_out_6_d23, arith_out_col_out_6_d24 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_6_q24 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_7, arith_out_col_out_7_d1, arith_out_col_out_7_d2, arith_out_col_out_7_d3, arith_out_col_out_7_d4, arith_out_col_out_7_d5, arith_out_col_out_7_d6, arith_out_col_out_7_d7, arith_out_col_out_7_d8, arith_out_col_out_7_d9, arith_out_col_out_7_d10, arith_out_col_out_7_d11, arith_out_col_out_7_d12, arith_out_col_out_7_d13, arith_out_col_out_7_d14, arith_out_col_out_7_d15, arith_out_col_out_7_d16, arith_out_col_out_7_d17, arith_out_col_out_7_d18, arith_out_col_out_7_d19, arith_out_col_out_7_d20, arith_out_col_out_7_d21, arith_out_col_out_7_d22, arith_out_col_out_7_d23 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_7_q23 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_8, arith_out_col_out_8_d1, arith_out_col_out_8_d2, arith_out_col_out_8_d3, arith_out_col_out_8_d4, arith_out_col_out_8_d5, arith_out_col_out_8_d6, arith_out_col_out_8_d7, arith_out_col_out_8_d8, arith_out_col_out_8_d9, arith_out_col_out_8_d10, arith_out_col_out_8_d11, arith_out_col_out_8_d12, arith_out_col_out_8_d13, arith_out_col_out_8_d14, arith_out_col_out_8_d15, arith_out_col_out_8_d16, arith_out_col_out_8_d17, arith_out_col_out_8_d18, arith_out_col_out_8_d19, arith_out_col_out_8_d20, arith_out_col_out_8_d21, arith_out_col_out_8_d22 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_8_q22 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_9, arith_out_col_out_9_d1, arith_out_col_out_9_d2, arith_out_col_out_9_d3, arith_out_col_out_9_d4, arith_out_col_out_9_d5, arith_out_col_out_9_d6, arith_out_col_out_9_d7, arith_out_col_out_9_d8, arith_out_col_out_9_d9, arith_out_col_out_9_d10, arith_out_col_out_9_d11, arith_out_col_out_9_d12, arith_out_col_out_9_d13, arith_out_col_out_9_d14, arith_out_col_out_9_d15, arith_out_col_out_9_d16, arith_out_col_out_9_d17, arith_out_col_out_9_d18, arith_out_col_out_9_d19, arith_out_col_out_9_d20, arith_out_col_out_9_d21 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_9_q21 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_10, arith_out_col_out_10_d1, arith_out_col_out_10_d2, arith_out_col_out_10_d3, arith_out_col_out_10_d4, arith_out_col_out_10_d5, arith_out_col_out_10_d6, arith_out_col_out_10_d7, arith_out_col_out_10_d8, arith_out_col_out_10_d9, arith_out_col_out_10_d10, arith_out_col_out_10_d11, arith_out_col_out_10_d12, arith_out_col_out_10_d13, arith_out_col_out_10_d14, arith_out_col_out_10_d15, arith_out_col_out_10_d16, arith_out_col_out_10_d17, arith_out_col_out_10_d18, arith_out_col_out_10_d19, arith_out_col_out_10_d20 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_10_q20 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_11, arith_out_col_out_11_d1, arith_out_col_out_11_d2, arith_out_col_out_11_d3, arith_out_col_out_11_d4, arith_out_col_out_11_d5, arith_out_col_out_11_d6, arith_out_col_out_11_d7, arith_out_col_out_11_d8, arith_out_col_out_11_d9, arith_out_col_out_11_d10, arith_out_col_out_11_d11, arith_out_col_out_11_d12, arith_out_col_out_11_d13, arith_out_col_out_11_d14, arith_out_col_out_11_d15, arith_out_col_out_11_d16, arith_out_col_out_11_d17, arith_out_col_out_11_d18, arith_out_col_out_11_d19 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_11_q19 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_12, arith_out_col_out_12_d1, arith_out_col_out_12_d2, arith_out_col_out_12_d3, arith_out_col_out_12_d4, arith_out_col_out_12_d5, arith_out_col_out_12_d6, arith_out_col_out_12_d7, arith_out_col_out_12_d8, arith_out_col_out_12_d9, arith_out_col_out_12_d10, arith_out_col_out_12_d11, arith_out_col_out_12_d12, arith_out_col_out_12_d13, arith_out_col_out_12_d14, arith_out_col_out_12_d15, arith_out_col_out_12_d16, arith_out_col_out_12_d17, arith_out_col_out_12_d18 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_12_q18 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_13, arith_out_col_out_13_d1, arith_out_col_out_13_d2, arith_out_col_out_13_d3, arith_out_col_out_13_d4, arith_out_col_out_13_d5, arith_out_col_out_13_d6, arith_out_col_out_13_d7, arith_out_col_out_13_d8, arith_out_col_out_13_d9, arith_out_col_out_13_d10, arith_out_col_out_13_d11, arith_out_col_out_13_d12, arith_out_col_out_13_d13, arith_out_col_out_13_d14, arith_out_col_out_13_d15, arith_out_col_out_13_d16, arith_out_col_out_13_d17 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_13_q17 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_14, arith_out_col_out_14_d1, arith_out_col_out_14_d2, arith_out_col_out_14_d3, arith_out_col_out_14_d4, arith_out_col_out_14_d5, arith_out_col_out_14_d6, arith_out_col_out_14_d7, arith_out_col_out_14_d8, arith_out_col_out_14_d9, arith_out_col_out_14_d10, arith_out_col_out_14_d11, arith_out_col_out_14_d12, arith_out_col_out_14_d13, arith_out_col_out_14_d14, arith_out_col_out_14_d15, arith_out_col_out_14_d16 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_14_q16 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_15, arith_out_col_out_15_d1, arith_out_col_out_15_d2, arith_out_col_out_15_d3, arith_out_col_out_15_d4, arith_out_col_out_15_d5, arith_out_col_out_15_d6, arith_out_col_out_15_d7, arith_out_col_out_15_d8, arith_out_col_out_15_d9, arith_out_col_out_15_d10, arith_out_col_out_15_d11, arith_out_col_out_15_d12, arith_out_col_out_15_d13, arith_out_col_out_15_d14, arith_out_col_out_15_d15 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_15_q15 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_16, arith_out_col_out_16_d1, arith_out_col_out_16_d2, arith_out_col_out_16_d3, arith_out_col_out_16_d4, arith_out_col_out_16_d5, arith_out_col_out_16_d6, arith_out_col_out_16_d7, arith_out_col_out_16_d8, arith_out_col_out_16_d9, arith_out_col_out_16_d10, arith_out_col_out_16_d11, arith_out_col_out_16_d12, arith_out_col_out_16_d13, arith_out_col_out_16_d14 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_16_q14 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_17, arith_out_col_out_17_d1, arith_out_col_out_17_d2, arith_out_col_out_17_d3, arith_out_col_out_17_d4, arith_out_col_out_17_d5, arith_out_col_out_17_d6, arith_out_col_out_17_d7, arith_out_col_out_17_d8, arith_out_col_out_17_d9, arith_out_col_out_17_d10, arith_out_col_out_17_d11, arith_out_col_out_17_d12, arith_out_col_out_17_d13 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_17_q13 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_18, arith_out_col_out_18_d1, arith_out_col_out_18_d2, arith_out_col_out_18_d3, arith_out_col_out_18_d4, arith_out_col_out_18_d5, arith_out_col_out_18_d6, arith_out_col_out_18_d7, arith_out_col_out_18_d8, arith_out_col_out_18_d9, arith_out_col_out_18_d10, arith_out_col_out_18_d11, arith_out_col_out_18_d12 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_18_q12 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_19, arith_out_col_out_19_d1, arith_out_col_out_19_d2, arith_out_col_out_19_d3, arith_out_col_out_19_d4, arith_out_col_out_19_d5, arith_out_col_out_19_d6, arith_out_col_out_19_d7, arith_out_col_out_19_d8, arith_out_col_out_19_d9, arith_out_col_out_19_d10, arith_out_col_out_19_d11 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_19_q11 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_20, arith_out_col_out_20_d1, arith_out_col_out_20_d2, arith_out_col_out_20_d3, arith_out_col_out_20_d4, arith_out_col_out_20_d5, arith_out_col_out_20_d6, arith_out_col_out_20_d7, arith_out_col_out_20_d8, arith_out_col_out_20_d9, arith_out_col_out_20_d10 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_20_q10 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_21, arith_out_col_out_21_d1, arith_out_col_out_21_d2, arith_out_col_out_21_d3, arith_out_col_out_21_d4, arith_out_col_out_21_d5, arith_out_col_out_21_d6, arith_out_col_out_21_d7, arith_out_col_out_21_d8, arith_out_col_out_21_d9 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_21_q9 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_22, arith_out_col_out_22_d1, arith_out_col_out_22_d2, arith_out_col_out_22_d3, arith_out_col_out_22_d4, arith_out_col_out_22_d5, arith_out_col_out_22_d6, arith_out_col_out_22_d7, arith_out_col_out_22_d8 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_22_q8 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_23, arith_out_col_out_23_d1, arith_out_col_out_23_d2, arith_out_col_out_23_d3, arith_out_col_out_23_d4, arith_out_col_out_23_d5, arith_out_col_out_23_d6, arith_out_col_out_23_d7 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_23_q7 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_24, arith_out_col_out_24_d1, arith_out_col_out_24_d2, arith_out_col_out_24_d3, arith_out_col_out_24_d4, arith_out_col_out_24_d5, arith_out_col_out_24_d6 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_24_q6 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_25, arith_out_col_out_25_d1, arith_out_col_out_25_d2, arith_out_col_out_25_d3, arith_out_col_out_25_d4, arith_out_col_out_25_d5 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_25_q5 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_26, arith_out_col_out_26_d1, arith_out_col_out_26_d2, arith_out_col_out_26_d3, arith_out_col_out_26_d4 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_26_q4 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_27, arith_out_col_out_27_d1, arith_out_col_out_27_d2, arith_out_col_out_27_d3 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_27_q3 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_28, arith_out_col_out_28_d1, arith_out_col_out_28_d2 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_28_q2 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_29, arith_out_col_out_29_d1 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_29_q1 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_30 :  std_logic_vector(3 downto 0);
signal arith_out_col_out_30_q0 :  std_logic_vector(3 downto 0);
signal rows_i_arith : array_N_dense;
signal rows_i_s3 :  std_logic_vector(223 downto 0);
signal cols_j_arith : array_M_dense;
signal cols_j_s3 :  std_logic_vector(216 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            arith_in_row_1_d1 <=  arith_in_row_1;
            arith_in_row_2_d1 <=  arith_in_row_2;
            arith_in_row_2_d2 <=  arith_in_row_2_d1;
            arith_in_row_3_d1 <=  arith_in_row_3;
            arith_in_row_3_d2 <=  arith_in_row_3_d1;
            arith_in_row_3_d3 <=  arith_in_row_3_d2;
            arith_in_row_4_d1 <=  arith_in_row_4;
            arith_in_row_4_d2 <=  arith_in_row_4_d1;
            arith_in_row_4_d3 <=  arith_in_row_4_d2;
            arith_in_row_4_d4 <=  arith_in_row_4_d3;
            arith_in_row_5_d1 <=  arith_in_row_5;
            arith_in_row_5_d2 <=  arith_in_row_5_d1;
            arith_in_row_5_d3 <=  arith_in_row_5_d2;
            arith_in_row_5_d4 <=  arith_in_row_5_d3;
            arith_in_row_5_d5 <=  arith_in_row_5_d4;
            arith_in_row_6_d1 <=  arith_in_row_6;
            arith_in_row_6_d2 <=  arith_in_row_6_d1;
            arith_in_row_6_d3 <=  arith_in_row_6_d2;
            arith_in_row_6_d4 <=  arith_in_row_6_d3;
            arith_in_row_6_d5 <=  arith_in_row_6_d4;
            arith_in_row_6_d6 <=  arith_in_row_6_d5;
            arith_in_row_7_d1 <=  arith_in_row_7;
            arith_in_row_7_d2 <=  arith_in_row_7_d1;
            arith_in_row_7_d3 <=  arith_in_row_7_d2;
            arith_in_row_7_d4 <=  arith_in_row_7_d3;
            arith_in_row_7_d5 <=  arith_in_row_7_d4;
            arith_in_row_7_d6 <=  arith_in_row_7_d5;
            arith_in_row_7_d7 <=  arith_in_row_7_d6;
            arith_in_row_8_d1 <=  arith_in_row_8;
            arith_in_row_8_d2 <=  arith_in_row_8_d1;
            arith_in_row_8_d3 <=  arith_in_row_8_d2;
            arith_in_row_8_d4 <=  arith_in_row_8_d3;
            arith_in_row_8_d5 <=  arith_in_row_8_d4;
            arith_in_row_8_d6 <=  arith_in_row_8_d5;
            arith_in_row_8_d7 <=  arith_in_row_8_d6;
            arith_in_row_8_d8 <=  arith_in_row_8_d7;
            arith_in_row_9_d1 <=  arith_in_row_9;
            arith_in_row_9_d2 <=  arith_in_row_9_d1;
            arith_in_row_9_d3 <=  arith_in_row_9_d2;
            arith_in_row_9_d4 <=  arith_in_row_9_d3;
            arith_in_row_9_d5 <=  arith_in_row_9_d4;
            arith_in_row_9_d6 <=  arith_in_row_9_d5;
            arith_in_row_9_d7 <=  arith_in_row_9_d6;
            arith_in_row_9_d8 <=  arith_in_row_9_d7;
            arith_in_row_9_d9 <=  arith_in_row_9_d8;
            arith_in_row_10_d1 <=  arith_in_row_10;
            arith_in_row_10_d2 <=  arith_in_row_10_d1;
            arith_in_row_10_d3 <=  arith_in_row_10_d2;
            arith_in_row_10_d4 <=  arith_in_row_10_d3;
            arith_in_row_10_d5 <=  arith_in_row_10_d4;
            arith_in_row_10_d6 <=  arith_in_row_10_d5;
            arith_in_row_10_d7 <=  arith_in_row_10_d6;
            arith_in_row_10_d8 <=  arith_in_row_10_d7;
            arith_in_row_10_d9 <=  arith_in_row_10_d8;
            arith_in_row_10_d10 <=  arith_in_row_10_d9;
            arith_in_row_11_d1 <=  arith_in_row_11;
            arith_in_row_11_d2 <=  arith_in_row_11_d1;
            arith_in_row_11_d3 <=  arith_in_row_11_d2;
            arith_in_row_11_d4 <=  arith_in_row_11_d3;
            arith_in_row_11_d5 <=  arith_in_row_11_d4;
            arith_in_row_11_d6 <=  arith_in_row_11_d5;
            arith_in_row_11_d7 <=  arith_in_row_11_d6;
            arith_in_row_11_d8 <=  arith_in_row_11_d7;
            arith_in_row_11_d9 <=  arith_in_row_11_d8;
            arith_in_row_11_d10 <=  arith_in_row_11_d9;
            arith_in_row_11_d11 <=  arith_in_row_11_d10;
            arith_in_row_12_d1 <=  arith_in_row_12;
            arith_in_row_12_d2 <=  arith_in_row_12_d1;
            arith_in_row_12_d3 <=  arith_in_row_12_d2;
            arith_in_row_12_d4 <=  arith_in_row_12_d3;
            arith_in_row_12_d5 <=  arith_in_row_12_d4;
            arith_in_row_12_d6 <=  arith_in_row_12_d5;
            arith_in_row_12_d7 <=  arith_in_row_12_d6;
            arith_in_row_12_d8 <=  arith_in_row_12_d7;
            arith_in_row_12_d9 <=  arith_in_row_12_d8;
            arith_in_row_12_d10 <=  arith_in_row_12_d9;
            arith_in_row_12_d11 <=  arith_in_row_12_d10;
            arith_in_row_12_d12 <=  arith_in_row_12_d11;
            arith_in_row_13_d1 <=  arith_in_row_13;
            arith_in_row_13_d2 <=  arith_in_row_13_d1;
            arith_in_row_13_d3 <=  arith_in_row_13_d2;
            arith_in_row_13_d4 <=  arith_in_row_13_d3;
            arith_in_row_13_d5 <=  arith_in_row_13_d4;
            arith_in_row_13_d6 <=  arith_in_row_13_d5;
            arith_in_row_13_d7 <=  arith_in_row_13_d6;
            arith_in_row_13_d8 <=  arith_in_row_13_d7;
            arith_in_row_13_d9 <=  arith_in_row_13_d8;
            arith_in_row_13_d10 <=  arith_in_row_13_d9;
            arith_in_row_13_d11 <=  arith_in_row_13_d10;
            arith_in_row_13_d12 <=  arith_in_row_13_d11;
            arith_in_row_13_d13 <=  arith_in_row_13_d12;
            arith_in_row_14_d1 <=  arith_in_row_14;
            arith_in_row_14_d2 <=  arith_in_row_14_d1;
            arith_in_row_14_d3 <=  arith_in_row_14_d2;
            arith_in_row_14_d4 <=  arith_in_row_14_d3;
            arith_in_row_14_d5 <=  arith_in_row_14_d4;
            arith_in_row_14_d6 <=  arith_in_row_14_d5;
            arith_in_row_14_d7 <=  arith_in_row_14_d6;
            arith_in_row_14_d8 <=  arith_in_row_14_d7;
            arith_in_row_14_d9 <=  arith_in_row_14_d8;
            arith_in_row_14_d10 <=  arith_in_row_14_d9;
            arith_in_row_14_d11 <=  arith_in_row_14_d10;
            arith_in_row_14_d12 <=  arith_in_row_14_d11;
            arith_in_row_14_d13 <=  arith_in_row_14_d12;
            arith_in_row_14_d14 <=  arith_in_row_14_d13;
            arith_in_row_15_d1 <=  arith_in_row_15;
            arith_in_row_15_d2 <=  arith_in_row_15_d1;
            arith_in_row_15_d3 <=  arith_in_row_15_d2;
            arith_in_row_15_d4 <=  arith_in_row_15_d3;
            arith_in_row_15_d5 <=  arith_in_row_15_d4;
            arith_in_row_15_d6 <=  arith_in_row_15_d5;
            arith_in_row_15_d7 <=  arith_in_row_15_d6;
            arith_in_row_15_d8 <=  arith_in_row_15_d7;
            arith_in_row_15_d9 <=  arith_in_row_15_d8;
            arith_in_row_15_d10 <=  arith_in_row_15_d9;
            arith_in_row_15_d11 <=  arith_in_row_15_d10;
            arith_in_row_15_d12 <=  arith_in_row_15_d11;
            arith_in_row_15_d13 <=  arith_in_row_15_d12;
            arith_in_row_15_d14 <=  arith_in_row_15_d13;
            arith_in_row_15_d15 <=  arith_in_row_15_d14;
            arith_in_row_16_d1 <=  arith_in_row_16;
            arith_in_row_16_d2 <=  arith_in_row_16_d1;
            arith_in_row_16_d3 <=  arith_in_row_16_d2;
            arith_in_row_16_d4 <=  arith_in_row_16_d3;
            arith_in_row_16_d5 <=  arith_in_row_16_d4;
            arith_in_row_16_d6 <=  arith_in_row_16_d5;
            arith_in_row_16_d7 <=  arith_in_row_16_d6;
            arith_in_row_16_d8 <=  arith_in_row_16_d7;
            arith_in_row_16_d9 <=  arith_in_row_16_d8;
            arith_in_row_16_d10 <=  arith_in_row_16_d9;
            arith_in_row_16_d11 <=  arith_in_row_16_d10;
            arith_in_row_16_d12 <=  arith_in_row_16_d11;
            arith_in_row_16_d13 <=  arith_in_row_16_d12;
            arith_in_row_16_d14 <=  arith_in_row_16_d13;
            arith_in_row_16_d15 <=  arith_in_row_16_d14;
            arith_in_row_16_d16 <=  arith_in_row_16_d15;
            arith_in_row_17_d1 <=  arith_in_row_17;
            arith_in_row_17_d2 <=  arith_in_row_17_d1;
            arith_in_row_17_d3 <=  arith_in_row_17_d2;
            arith_in_row_17_d4 <=  arith_in_row_17_d3;
            arith_in_row_17_d5 <=  arith_in_row_17_d4;
            arith_in_row_17_d6 <=  arith_in_row_17_d5;
            arith_in_row_17_d7 <=  arith_in_row_17_d6;
            arith_in_row_17_d8 <=  arith_in_row_17_d7;
            arith_in_row_17_d9 <=  arith_in_row_17_d8;
            arith_in_row_17_d10 <=  arith_in_row_17_d9;
            arith_in_row_17_d11 <=  arith_in_row_17_d10;
            arith_in_row_17_d12 <=  arith_in_row_17_d11;
            arith_in_row_17_d13 <=  arith_in_row_17_d12;
            arith_in_row_17_d14 <=  arith_in_row_17_d13;
            arith_in_row_17_d15 <=  arith_in_row_17_d14;
            arith_in_row_17_d16 <=  arith_in_row_17_d15;
            arith_in_row_17_d17 <=  arith_in_row_17_d16;
            arith_in_row_18_d1 <=  arith_in_row_18;
            arith_in_row_18_d2 <=  arith_in_row_18_d1;
            arith_in_row_18_d3 <=  arith_in_row_18_d2;
            arith_in_row_18_d4 <=  arith_in_row_18_d3;
            arith_in_row_18_d5 <=  arith_in_row_18_d4;
            arith_in_row_18_d6 <=  arith_in_row_18_d5;
            arith_in_row_18_d7 <=  arith_in_row_18_d6;
            arith_in_row_18_d8 <=  arith_in_row_18_d7;
            arith_in_row_18_d9 <=  arith_in_row_18_d8;
            arith_in_row_18_d10 <=  arith_in_row_18_d9;
            arith_in_row_18_d11 <=  arith_in_row_18_d10;
            arith_in_row_18_d12 <=  arith_in_row_18_d11;
            arith_in_row_18_d13 <=  arith_in_row_18_d12;
            arith_in_row_18_d14 <=  arith_in_row_18_d13;
            arith_in_row_18_d15 <=  arith_in_row_18_d14;
            arith_in_row_18_d16 <=  arith_in_row_18_d15;
            arith_in_row_18_d17 <=  arith_in_row_18_d16;
            arith_in_row_18_d18 <=  arith_in_row_18_d17;
            arith_in_row_19_d1 <=  arith_in_row_19;
            arith_in_row_19_d2 <=  arith_in_row_19_d1;
            arith_in_row_19_d3 <=  arith_in_row_19_d2;
            arith_in_row_19_d4 <=  arith_in_row_19_d3;
            arith_in_row_19_d5 <=  arith_in_row_19_d4;
            arith_in_row_19_d6 <=  arith_in_row_19_d5;
            arith_in_row_19_d7 <=  arith_in_row_19_d6;
            arith_in_row_19_d8 <=  arith_in_row_19_d7;
            arith_in_row_19_d9 <=  arith_in_row_19_d8;
            arith_in_row_19_d10 <=  arith_in_row_19_d9;
            arith_in_row_19_d11 <=  arith_in_row_19_d10;
            arith_in_row_19_d12 <=  arith_in_row_19_d11;
            arith_in_row_19_d13 <=  arith_in_row_19_d12;
            arith_in_row_19_d14 <=  arith_in_row_19_d13;
            arith_in_row_19_d15 <=  arith_in_row_19_d14;
            arith_in_row_19_d16 <=  arith_in_row_19_d15;
            arith_in_row_19_d17 <=  arith_in_row_19_d16;
            arith_in_row_19_d18 <=  arith_in_row_19_d17;
            arith_in_row_19_d19 <=  arith_in_row_19_d18;
            arith_in_row_20_d1 <=  arith_in_row_20;
            arith_in_row_20_d2 <=  arith_in_row_20_d1;
            arith_in_row_20_d3 <=  arith_in_row_20_d2;
            arith_in_row_20_d4 <=  arith_in_row_20_d3;
            arith_in_row_20_d5 <=  arith_in_row_20_d4;
            arith_in_row_20_d6 <=  arith_in_row_20_d5;
            arith_in_row_20_d7 <=  arith_in_row_20_d6;
            arith_in_row_20_d8 <=  arith_in_row_20_d7;
            arith_in_row_20_d9 <=  arith_in_row_20_d8;
            arith_in_row_20_d10 <=  arith_in_row_20_d9;
            arith_in_row_20_d11 <=  arith_in_row_20_d10;
            arith_in_row_20_d12 <=  arith_in_row_20_d11;
            arith_in_row_20_d13 <=  arith_in_row_20_d12;
            arith_in_row_20_d14 <=  arith_in_row_20_d13;
            arith_in_row_20_d15 <=  arith_in_row_20_d14;
            arith_in_row_20_d16 <=  arith_in_row_20_d15;
            arith_in_row_20_d17 <=  arith_in_row_20_d16;
            arith_in_row_20_d18 <=  arith_in_row_20_d17;
            arith_in_row_20_d19 <=  arith_in_row_20_d18;
            arith_in_row_20_d20 <=  arith_in_row_20_d19;
            arith_in_row_21_d1 <=  arith_in_row_21;
            arith_in_row_21_d2 <=  arith_in_row_21_d1;
            arith_in_row_21_d3 <=  arith_in_row_21_d2;
            arith_in_row_21_d4 <=  arith_in_row_21_d3;
            arith_in_row_21_d5 <=  arith_in_row_21_d4;
            arith_in_row_21_d6 <=  arith_in_row_21_d5;
            arith_in_row_21_d7 <=  arith_in_row_21_d6;
            arith_in_row_21_d8 <=  arith_in_row_21_d7;
            arith_in_row_21_d9 <=  arith_in_row_21_d8;
            arith_in_row_21_d10 <=  arith_in_row_21_d9;
            arith_in_row_21_d11 <=  arith_in_row_21_d10;
            arith_in_row_21_d12 <=  arith_in_row_21_d11;
            arith_in_row_21_d13 <=  arith_in_row_21_d12;
            arith_in_row_21_d14 <=  arith_in_row_21_d13;
            arith_in_row_21_d15 <=  arith_in_row_21_d14;
            arith_in_row_21_d16 <=  arith_in_row_21_d15;
            arith_in_row_21_d17 <=  arith_in_row_21_d16;
            arith_in_row_21_d18 <=  arith_in_row_21_d17;
            arith_in_row_21_d19 <=  arith_in_row_21_d18;
            arith_in_row_21_d20 <=  arith_in_row_21_d19;
            arith_in_row_21_d21 <=  arith_in_row_21_d20;
            arith_in_row_22_d1 <=  arith_in_row_22;
            arith_in_row_22_d2 <=  arith_in_row_22_d1;
            arith_in_row_22_d3 <=  arith_in_row_22_d2;
            arith_in_row_22_d4 <=  arith_in_row_22_d3;
            arith_in_row_22_d5 <=  arith_in_row_22_d4;
            arith_in_row_22_d6 <=  arith_in_row_22_d5;
            arith_in_row_22_d7 <=  arith_in_row_22_d6;
            arith_in_row_22_d8 <=  arith_in_row_22_d7;
            arith_in_row_22_d9 <=  arith_in_row_22_d8;
            arith_in_row_22_d10 <=  arith_in_row_22_d9;
            arith_in_row_22_d11 <=  arith_in_row_22_d10;
            arith_in_row_22_d12 <=  arith_in_row_22_d11;
            arith_in_row_22_d13 <=  arith_in_row_22_d12;
            arith_in_row_22_d14 <=  arith_in_row_22_d13;
            arith_in_row_22_d15 <=  arith_in_row_22_d14;
            arith_in_row_22_d16 <=  arith_in_row_22_d15;
            arith_in_row_22_d17 <=  arith_in_row_22_d16;
            arith_in_row_22_d18 <=  arith_in_row_22_d17;
            arith_in_row_22_d19 <=  arith_in_row_22_d18;
            arith_in_row_22_d20 <=  arith_in_row_22_d19;
            arith_in_row_22_d21 <=  arith_in_row_22_d20;
            arith_in_row_22_d22 <=  arith_in_row_22_d21;
            arith_in_row_23_d1 <=  arith_in_row_23;
            arith_in_row_23_d2 <=  arith_in_row_23_d1;
            arith_in_row_23_d3 <=  arith_in_row_23_d2;
            arith_in_row_23_d4 <=  arith_in_row_23_d3;
            arith_in_row_23_d5 <=  arith_in_row_23_d4;
            arith_in_row_23_d6 <=  arith_in_row_23_d5;
            arith_in_row_23_d7 <=  arith_in_row_23_d6;
            arith_in_row_23_d8 <=  arith_in_row_23_d7;
            arith_in_row_23_d9 <=  arith_in_row_23_d8;
            arith_in_row_23_d10 <=  arith_in_row_23_d9;
            arith_in_row_23_d11 <=  arith_in_row_23_d10;
            arith_in_row_23_d12 <=  arith_in_row_23_d11;
            arith_in_row_23_d13 <=  arith_in_row_23_d12;
            arith_in_row_23_d14 <=  arith_in_row_23_d13;
            arith_in_row_23_d15 <=  arith_in_row_23_d14;
            arith_in_row_23_d16 <=  arith_in_row_23_d15;
            arith_in_row_23_d17 <=  arith_in_row_23_d16;
            arith_in_row_23_d18 <=  arith_in_row_23_d17;
            arith_in_row_23_d19 <=  arith_in_row_23_d18;
            arith_in_row_23_d20 <=  arith_in_row_23_d19;
            arith_in_row_23_d21 <=  arith_in_row_23_d20;
            arith_in_row_23_d22 <=  arith_in_row_23_d21;
            arith_in_row_23_d23 <=  arith_in_row_23_d22;
            arith_in_row_24_d1 <=  arith_in_row_24;
            arith_in_row_24_d2 <=  arith_in_row_24_d1;
            arith_in_row_24_d3 <=  arith_in_row_24_d2;
            arith_in_row_24_d4 <=  arith_in_row_24_d3;
            arith_in_row_24_d5 <=  arith_in_row_24_d4;
            arith_in_row_24_d6 <=  arith_in_row_24_d5;
            arith_in_row_24_d7 <=  arith_in_row_24_d6;
            arith_in_row_24_d8 <=  arith_in_row_24_d7;
            arith_in_row_24_d9 <=  arith_in_row_24_d8;
            arith_in_row_24_d10 <=  arith_in_row_24_d9;
            arith_in_row_24_d11 <=  arith_in_row_24_d10;
            arith_in_row_24_d12 <=  arith_in_row_24_d11;
            arith_in_row_24_d13 <=  arith_in_row_24_d12;
            arith_in_row_24_d14 <=  arith_in_row_24_d13;
            arith_in_row_24_d15 <=  arith_in_row_24_d14;
            arith_in_row_24_d16 <=  arith_in_row_24_d15;
            arith_in_row_24_d17 <=  arith_in_row_24_d16;
            arith_in_row_24_d18 <=  arith_in_row_24_d17;
            arith_in_row_24_d19 <=  arith_in_row_24_d18;
            arith_in_row_24_d20 <=  arith_in_row_24_d19;
            arith_in_row_24_d21 <=  arith_in_row_24_d20;
            arith_in_row_24_d22 <=  arith_in_row_24_d21;
            arith_in_row_24_d23 <=  arith_in_row_24_d22;
            arith_in_row_24_d24 <=  arith_in_row_24_d23;
            arith_in_row_25_d1 <=  arith_in_row_25;
            arith_in_row_25_d2 <=  arith_in_row_25_d1;
            arith_in_row_25_d3 <=  arith_in_row_25_d2;
            arith_in_row_25_d4 <=  arith_in_row_25_d3;
            arith_in_row_25_d5 <=  arith_in_row_25_d4;
            arith_in_row_25_d6 <=  arith_in_row_25_d5;
            arith_in_row_25_d7 <=  arith_in_row_25_d6;
            arith_in_row_25_d8 <=  arith_in_row_25_d7;
            arith_in_row_25_d9 <=  arith_in_row_25_d8;
            arith_in_row_25_d10 <=  arith_in_row_25_d9;
            arith_in_row_25_d11 <=  arith_in_row_25_d10;
            arith_in_row_25_d12 <=  arith_in_row_25_d11;
            arith_in_row_25_d13 <=  arith_in_row_25_d12;
            arith_in_row_25_d14 <=  arith_in_row_25_d13;
            arith_in_row_25_d15 <=  arith_in_row_25_d14;
            arith_in_row_25_d16 <=  arith_in_row_25_d15;
            arith_in_row_25_d17 <=  arith_in_row_25_d16;
            arith_in_row_25_d18 <=  arith_in_row_25_d17;
            arith_in_row_25_d19 <=  arith_in_row_25_d18;
            arith_in_row_25_d20 <=  arith_in_row_25_d19;
            arith_in_row_25_d21 <=  arith_in_row_25_d20;
            arith_in_row_25_d22 <=  arith_in_row_25_d21;
            arith_in_row_25_d23 <=  arith_in_row_25_d22;
            arith_in_row_25_d24 <=  arith_in_row_25_d23;
            arith_in_row_25_d25 <=  arith_in_row_25_d24;
            arith_in_row_26_d1 <=  arith_in_row_26;
            arith_in_row_26_d2 <=  arith_in_row_26_d1;
            arith_in_row_26_d3 <=  arith_in_row_26_d2;
            arith_in_row_26_d4 <=  arith_in_row_26_d3;
            arith_in_row_26_d5 <=  arith_in_row_26_d4;
            arith_in_row_26_d6 <=  arith_in_row_26_d5;
            arith_in_row_26_d7 <=  arith_in_row_26_d6;
            arith_in_row_26_d8 <=  arith_in_row_26_d7;
            arith_in_row_26_d9 <=  arith_in_row_26_d8;
            arith_in_row_26_d10 <=  arith_in_row_26_d9;
            arith_in_row_26_d11 <=  arith_in_row_26_d10;
            arith_in_row_26_d12 <=  arith_in_row_26_d11;
            arith_in_row_26_d13 <=  arith_in_row_26_d12;
            arith_in_row_26_d14 <=  arith_in_row_26_d13;
            arith_in_row_26_d15 <=  arith_in_row_26_d14;
            arith_in_row_26_d16 <=  arith_in_row_26_d15;
            arith_in_row_26_d17 <=  arith_in_row_26_d16;
            arith_in_row_26_d18 <=  arith_in_row_26_d17;
            arith_in_row_26_d19 <=  arith_in_row_26_d18;
            arith_in_row_26_d20 <=  arith_in_row_26_d19;
            arith_in_row_26_d21 <=  arith_in_row_26_d20;
            arith_in_row_26_d22 <=  arith_in_row_26_d21;
            arith_in_row_26_d23 <=  arith_in_row_26_d22;
            arith_in_row_26_d24 <=  arith_in_row_26_d23;
            arith_in_row_26_d25 <=  arith_in_row_26_d24;
            arith_in_row_26_d26 <=  arith_in_row_26_d25;
            arith_in_row_27_d1 <=  arith_in_row_27;
            arith_in_row_27_d2 <=  arith_in_row_27_d1;
            arith_in_row_27_d3 <=  arith_in_row_27_d2;
            arith_in_row_27_d4 <=  arith_in_row_27_d3;
            arith_in_row_27_d5 <=  arith_in_row_27_d4;
            arith_in_row_27_d6 <=  arith_in_row_27_d5;
            arith_in_row_27_d7 <=  arith_in_row_27_d6;
            arith_in_row_27_d8 <=  arith_in_row_27_d7;
            arith_in_row_27_d9 <=  arith_in_row_27_d8;
            arith_in_row_27_d10 <=  arith_in_row_27_d9;
            arith_in_row_27_d11 <=  arith_in_row_27_d10;
            arith_in_row_27_d12 <=  arith_in_row_27_d11;
            arith_in_row_27_d13 <=  arith_in_row_27_d12;
            arith_in_row_27_d14 <=  arith_in_row_27_d13;
            arith_in_row_27_d15 <=  arith_in_row_27_d14;
            arith_in_row_27_d16 <=  arith_in_row_27_d15;
            arith_in_row_27_d17 <=  arith_in_row_27_d16;
            arith_in_row_27_d18 <=  arith_in_row_27_d17;
            arith_in_row_27_d19 <=  arith_in_row_27_d18;
            arith_in_row_27_d20 <=  arith_in_row_27_d19;
            arith_in_row_27_d21 <=  arith_in_row_27_d20;
            arith_in_row_27_d22 <=  arith_in_row_27_d21;
            arith_in_row_27_d23 <=  arith_in_row_27_d22;
            arith_in_row_27_d24 <=  arith_in_row_27_d23;
            arith_in_row_27_d25 <=  arith_in_row_27_d24;
            arith_in_row_27_d26 <=  arith_in_row_27_d25;
            arith_in_row_27_d27 <=  arith_in_row_27_d26;
            arith_in_row_28_d1 <=  arith_in_row_28;
            arith_in_row_28_d2 <=  arith_in_row_28_d1;
            arith_in_row_28_d3 <=  arith_in_row_28_d2;
            arith_in_row_28_d4 <=  arith_in_row_28_d3;
            arith_in_row_28_d5 <=  arith_in_row_28_d4;
            arith_in_row_28_d6 <=  arith_in_row_28_d5;
            arith_in_row_28_d7 <=  arith_in_row_28_d6;
            arith_in_row_28_d8 <=  arith_in_row_28_d7;
            arith_in_row_28_d9 <=  arith_in_row_28_d8;
            arith_in_row_28_d10 <=  arith_in_row_28_d9;
            arith_in_row_28_d11 <=  arith_in_row_28_d10;
            arith_in_row_28_d12 <=  arith_in_row_28_d11;
            arith_in_row_28_d13 <=  arith_in_row_28_d12;
            arith_in_row_28_d14 <=  arith_in_row_28_d13;
            arith_in_row_28_d15 <=  arith_in_row_28_d14;
            arith_in_row_28_d16 <=  arith_in_row_28_d15;
            arith_in_row_28_d17 <=  arith_in_row_28_d16;
            arith_in_row_28_d18 <=  arith_in_row_28_d17;
            arith_in_row_28_d19 <=  arith_in_row_28_d18;
            arith_in_row_28_d20 <=  arith_in_row_28_d19;
            arith_in_row_28_d21 <=  arith_in_row_28_d20;
            arith_in_row_28_d22 <=  arith_in_row_28_d21;
            arith_in_row_28_d23 <=  arith_in_row_28_d22;
            arith_in_row_28_d24 <=  arith_in_row_28_d23;
            arith_in_row_28_d25 <=  arith_in_row_28_d24;
            arith_in_row_28_d26 <=  arith_in_row_28_d25;
            arith_in_row_28_d27 <=  arith_in_row_28_d26;
            arith_in_row_28_d28 <=  arith_in_row_28_d27;
            arith_in_row_29_d1 <=  arith_in_row_29;
            arith_in_row_29_d2 <=  arith_in_row_29_d1;
            arith_in_row_29_d3 <=  arith_in_row_29_d2;
            arith_in_row_29_d4 <=  arith_in_row_29_d3;
            arith_in_row_29_d5 <=  arith_in_row_29_d4;
            arith_in_row_29_d6 <=  arith_in_row_29_d5;
            arith_in_row_29_d7 <=  arith_in_row_29_d6;
            arith_in_row_29_d8 <=  arith_in_row_29_d7;
            arith_in_row_29_d9 <=  arith_in_row_29_d8;
            arith_in_row_29_d10 <=  arith_in_row_29_d9;
            arith_in_row_29_d11 <=  arith_in_row_29_d10;
            arith_in_row_29_d12 <=  arith_in_row_29_d11;
            arith_in_row_29_d13 <=  arith_in_row_29_d12;
            arith_in_row_29_d14 <=  arith_in_row_29_d13;
            arith_in_row_29_d15 <=  arith_in_row_29_d14;
            arith_in_row_29_d16 <=  arith_in_row_29_d15;
            arith_in_row_29_d17 <=  arith_in_row_29_d16;
            arith_in_row_29_d18 <=  arith_in_row_29_d17;
            arith_in_row_29_d19 <=  arith_in_row_29_d18;
            arith_in_row_29_d20 <=  arith_in_row_29_d19;
            arith_in_row_29_d21 <=  arith_in_row_29_d20;
            arith_in_row_29_d22 <=  arith_in_row_29_d21;
            arith_in_row_29_d23 <=  arith_in_row_29_d22;
            arith_in_row_29_d24 <=  arith_in_row_29_d23;
            arith_in_row_29_d25 <=  arith_in_row_29_d24;
            arith_in_row_29_d26 <=  arith_in_row_29_d25;
            arith_in_row_29_d27 <=  arith_in_row_29_d26;
            arith_in_row_29_d28 <=  arith_in_row_29_d27;
            arith_in_row_29_d29 <=  arith_in_row_29_d28;
            arith_in_row_30_d1 <=  arith_in_row_30;
            arith_in_row_30_d2 <=  arith_in_row_30_d1;
            arith_in_row_30_d3 <=  arith_in_row_30_d2;
            arith_in_row_30_d4 <=  arith_in_row_30_d3;
            arith_in_row_30_d5 <=  arith_in_row_30_d4;
            arith_in_row_30_d6 <=  arith_in_row_30_d5;
            arith_in_row_30_d7 <=  arith_in_row_30_d6;
            arith_in_row_30_d8 <=  arith_in_row_30_d7;
            arith_in_row_30_d9 <=  arith_in_row_30_d8;
            arith_in_row_30_d10 <=  arith_in_row_30_d9;
            arith_in_row_30_d11 <=  arith_in_row_30_d10;
            arith_in_row_30_d12 <=  arith_in_row_30_d11;
            arith_in_row_30_d13 <=  arith_in_row_30_d12;
            arith_in_row_30_d14 <=  arith_in_row_30_d13;
            arith_in_row_30_d15 <=  arith_in_row_30_d14;
            arith_in_row_30_d16 <=  arith_in_row_30_d15;
            arith_in_row_30_d17 <=  arith_in_row_30_d16;
            arith_in_row_30_d18 <=  arith_in_row_30_d17;
            arith_in_row_30_d19 <=  arith_in_row_30_d18;
            arith_in_row_30_d20 <=  arith_in_row_30_d19;
            arith_in_row_30_d21 <=  arith_in_row_30_d20;
            arith_in_row_30_d22 <=  arith_in_row_30_d21;
            arith_in_row_30_d23 <=  arith_in_row_30_d22;
            arith_in_row_30_d24 <=  arith_in_row_30_d23;
            arith_in_row_30_d25 <=  arith_in_row_30_d24;
            arith_in_row_30_d26 <=  arith_in_row_30_d25;
            arith_in_row_30_d27 <=  arith_in_row_30_d26;
            arith_in_row_30_d28 <=  arith_in_row_30_d27;
            arith_in_row_30_d29 <=  arith_in_row_30_d28;
            arith_in_row_30_d30 <=  arith_in_row_30_d29;
            arith_in_row_31_d1 <=  arith_in_row_31;
            arith_in_row_31_d2 <=  arith_in_row_31_d1;
            arith_in_row_31_d3 <=  arith_in_row_31_d2;
            arith_in_row_31_d4 <=  arith_in_row_31_d3;
            arith_in_row_31_d5 <=  arith_in_row_31_d4;
            arith_in_row_31_d6 <=  arith_in_row_31_d5;
            arith_in_row_31_d7 <=  arith_in_row_31_d6;
            arith_in_row_31_d8 <=  arith_in_row_31_d7;
            arith_in_row_31_d9 <=  arith_in_row_31_d8;
            arith_in_row_31_d10 <=  arith_in_row_31_d9;
            arith_in_row_31_d11 <=  arith_in_row_31_d10;
            arith_in_row_31_d12 <=  arith_in_row_31_d11;
            arith_in_row_31_d13 <=  arith_in_row_31_d12;
            arith_in_row_31_d14 <=  arith_in_row_31_d13;
            arith_in_row_31_d15 <=  arith_in_row_31_d14;
            arith_in_row_31_d16 <=  arith_in_row_31_d15;
            arith_in_row_31_d17 <=  arith_in_row_31_d16;
            arith_in_row_31_d18 <=  arith_in_row_31_d17;
            arith_in_row_31_d19 <=  arith_in_row_31_d18;
            arith_in_row_31_d20 <=  arith_in_row_31_d19;
            arith_in_row_31_d21 <=  arith_in_row_31_d20;
            arith_in_row_31_d22 <=  arith_in_row_31_d21;
            arith_in_row_31_d23 <=  arith_in_row_31_d22;
            arith_in_row_31_d24 <=  arith_in_row_31_d23;
            arith_in_row_31_d25 <=  arith_in_row_31_d24;
            arith_in_row_31_d26 <=  arith_in_row_31_d25;
            arith_in_row_31_d27 <=  arith_in_row_31_d26;
            arith_in_row_31_d28 <=  arith_in_row_31_d27;
            arith_in_row_31_d29 <=  arith_in_row_31_d28;
            arith_in_row_31_d30 <=  arith_in_row_31_d29;
            arith_in_row_31_d31 <=  arith_in_row_31_d30;
            arith_in_col_1_d1 <=  arith_in_col_1;
            arith_in_col_2_d1 <=  arith_in_col_2;
            arith_in_col_2_d2 <=  arith_in_col_2_d1;
            arith_in_col_3_d1 <=  arith_in_col_3;
            arith_in_col_3_d2 <=  arith_in_col_3_d1;
            arith_in_col_3_d3 <=  arith_in_col_3_d2;
            arith_in_col_4_d1 <=  arith_in_col_4;
            arith_in_col_4_d2 <=  arith_in_col_4_d1;
            arith_in_col_4_d3 <=  arith_in_col_4_d2;
            arith_in_col_4_d4 <=  arith_in_col_4_d3;
            arith_in_col_5_d1 <=  arith_in_col_5;
            arith_in_col_5_d2 <=  arith_in_col_5_d1;
            arith_in_col_5_d3 <=  arith_in_col_5_d2;
            arith_in_col_5_d4 <=  arith_in_col_5_d3;
            arith_in_col_5_d5 <=  arith_in_col_5_d4;
            arith_in_col_6_d1 <=  arith_in_col_6;
            arith_in_col_6_d2 <=  arith_in_col_6_d1;
            arith_in_col_6_d3 <=  arith_in_col_6_d2;
            arith_in_col_6_d4 <=  arith_in_col_6_d3;
            arith_in_col_6_d5 <=  arith_in_col_6_d4;
            arith_in_col_6_d6 <=  arith_in_col_6_d5;
            arith_in_col_7_d1 <=  arith_in_col_7;
            arith_in_col_7_d2 <=  arith_in_col_7_d1;
            arith_in_col_7_d3 <=  arith_in_col_7_d2;
            arith_in_col_7_d4 <=  arith_in_col_7_d3;
            arith_in_col_7_d5 <=  arith_in_col_7_d4;
            arith_in_col_7_d6 <=  arith_in_col_7_d5;
            arith_in_col_7_d7 <=  arith_in_col_7_d6;
            arith_in_col_8_d1 <=  arith_in_col_8;
            arith_in_col_8_d2 <=  arith_in_col_8_d1;
            arith_in_col_8_d3 <=  arith_in_col_8_d2;
            arith_in_col_8_d4 <=  arith_in_col_8_d3;
            arith_in_col_8_d5 <=  arith_in_col_8_d4;
            arith_in_col_8_d6 <=  arith_in_col_8_d5;
            arith_in_col_8_d7 <=  arith_in_col_8_d6;
            arith_in_col_8_d8 <=  arith_in_col_8_d7;
            arith_in_col_9_d1 <=  arith_in_col_9;
            arith_in_col_9_d2 <=  arith_in_col_9_d1;
            arith_in_col_9_d3 <=  arith_in_col_9_d2;
            arith_in_col_9_d4 <=  arith_in_col_9_d3;
            arith_in_col_9_d5 <=  arith_in_col_9_d4;
            arith_in_col_9_d6 <=  arith_in_col_9_d5;
            arith_in_col_9_d7 <=  arith_in_col_9_d6;
            arith_in_col_9_d8 <=  arith_in_col_9_d7;
            arith_in_col_9_d9 <=  arith_in_col_9_d8;
            arith_in_col_10_d1 <=  arith_in_col_10;
            arith_in_col_10_d2 <=  arith_in_col_10_d1;
            arith_in_col_10_d3 <=  arith_in_col_10_d2;
            arith_in_col_10_d4 <=  arith_in_col_10_d3;
            arith_in_col_10_d5 <=  arith_in_col_10_d4;
            arith_in_col_10_d6 <=  arith_in_col_10_d5;
            arith_in_col_10_d7 <=  arith_in_col_10_d6;
            arith_in_col_10_d8 <=  arith_in_col_10_d7;
            arith_in_col_10_d9 <=  arith_in_col_10_d8;
            arith_in_col_10_d10 <=  arith_in_col_10_d9;
            arith_in_col_11_d1 <=  arith_in_col_11;
            arith_in_col_11_d2 <=  arith_in_col_11_d1;
            arith_in_col_11_d3 <=  arith_in_col_11_d2;
            arith_in_col_11_d4 <=  arith_in_col_11_d3;
            arith_in_col_11_d5 <=  arith_in_col_11_d4;
            arith_in_col_11_d6 <=  arith_in_col_11_d5;
            arith_in_col_11_d7 <=  arith_in_col_11_d6;
            arith_in_col_11_d8 <=  arith_in_col_11_d7;
            arith_in_col_11_d9 <=  arith_in_col_11_d8;
            arith_in_col_11_d10 <=  arith_in_col_11_d9;
            arith_in_col_11_d11 <=  arith_in_col_11_d10;
            arith_in_col_12_d1 <=  arith_in_col_12;
            arith_in_col_12_d2 <=  arith_in_col_12_d1;
            arith_in_col_12_d3 <=  arith_in_col_12_d2;
            arith_in_col_12_d4 <=  arith_in_col_12_d3;
            arith_in_col_12_d5 <=  arith_in_col_12_d4;
            arith_in_col_12_d6 <=  arith_in_col_12_d5;
            arith_in_col_12_d7 <=  arith_in_col_12_d6;
            arith_in_col_12_d8 <=  arith_in_col_12_d7;
            arith_in_col_12_d9 <=  arith_in_col_12_d8;
            arith_in_col_12_d10 <=  arith_in_col_12_d9;
            arith_in_col_12_d11 <=  arith_in_col_12_d10;
            arith_in_col_12_d12 <=  arith_in_col_12_d11;
            arith_in_col_13_d1 <=  arith_in_col_13;
            arith_in_col_13_d2 <=  arith_in_col_13_d1;
            arith_in_col_13_d3 <=  arith_in_col_13_d2;
            arith_in_col_13_d4 <=  arith_in_col_13_d3;
            arith_in_col_13_d5 <=  arith_in_col_13_d4;
            arith_in_col_13_d6 <=  arith_in_col_13_d5;
            arith_in_col_13_d7 <=  arith_in_col_13_d6;
            arith_in_col_13_d8 <=  arith_in_col_13_d7;
            arith_in_col_13_d9 <=  arith_in_col_13_d8;
            arith_in_col_13_d10 <=  arith_in_col_13_d9;
            arith_in_col_13_d11 <=  arith_in_col_13_d10;
            arith_in_col_13_d12 <=  arith_in_col_13_d11;
            arith_in_col_13_d13 <=  arith_in_col_13_d12;
            arith_in_col_14_d1 <=  arith_in_col_14;
            arith_in_col_14_d2 <=  arith_in_col_14_d1;
            arith_in_col_14_d3 <=  arith_in_col_14_d2;
            arith_in_col_14_d4 <=  arith_in_col_14_d3;
            arith_in_col_14_d5 <=  arith_in_col_14_d4;
            arith_in_col_14_d6 <=  arith_in_col_14_d5;
            arith_in_col_14_d7 <=  arith_in_col_14_d6;
            arith_in_col_14_d8 <=  arith_in_col_14_d7;
            arith_in_col_14_d9 <=  arith_in_col_14_d8;
            arith_in_col_14_d10 <=  arith_in_col_14_d9;
            arith_in_col_14_d11 <=  arith_in_col_14_d10;
            arith_in_col_14_d12 <=  arith_in_col_14_d11;
            arith_in_col_14_d13 <=  arith_in_col_14_d12;
            arith_in_col_14_d14 <=  arith_in_col_14_d13;
            arith_in_col_15_d1 <=  arith_in_col_15;
            arith_in_col_15_d2 <=  arith_in_col_15_d1;
            arith_in_col_15_d3 <=  arith_in_col_15_d2;
            arith_in_col_15_d4 <=  arith_in_col_15_d3;
            arith_in_col_15_d5 <=  arith_in_col_15_d4;
            arith_in_col_15_d6 <=  arith_in_col_15_d5;
            arith_in_col_15_d7 <=  arith_in_col_15_d6;
            arith_in_col_15_d8 <=  arith_in_col_15_d7;
            arith_in_col_15_d9 <=  arith_in_col_15_d8;
            arith_in_col_15_d10 <=  arith_in_col_15_d9;
            arith_in_col_15_d11 <=  arith_in_col_15_d10;
            arith_in_col_15_d12 <=  arith_in_col_15_d11;
            arith_in_col_15_d13 <=  arith_in_col_15_d12;
            arith_in_col_15_d14 <=  arith_in_col_15_d13;
            arith_in_col_15_d15 <=  arith_in_col_15_d14;
            arith_in_col_16_d1 <=  arith_in_col_16;
            arith_in_col_16_d2 <=  arith_in_col_16_d1;
            arith_in_col_16_d3 <=  arith_in_col_16_d2;
            arith_in_col_16_d4 <=  arith_in_col_16_d3;
            arith_in_col_16_d5 <=  arith_in_col_16_d4;
            arith_in_col_16_d6 <=  arith_in_col_16_d5;
            arith_in_col_16_d7 <=  arith_in_col_16_d6;
            arith_in_col_16_d8 <=  arith_in_col_16_d7;
            arith_in_col_16_d9 <=  arith_in_col_16_d8;
            arith_in_col_16_d10 <=  arith_in_col_16_d9;
            arith_in_col_16_d11 <=  arith_in_col_16_d10;
            arith_in_col_16_d12 <=  arith_in_col_16_d11;
            arith_in_col_16_d13 <=  arith_in_col_16_d12;
            arith_in_col_16_d14 <=  arith_in_col_16_d13;
            arith_in_col_16_d15 <=  arith_in_col_16_d14;
            arith_in_col_16_d16 <=  arith_in_col_16_d15;
            arith_in_col_17_d1 <=  arith_in_col_17;
            arith_in_col_17_d2 <=  arith_in_col_17_d1;
            arith_in_col_17_d3 <=  arith_in_col_17_d2;
            arith_in_col_17_d4 <=  arith_in_col_17_d3;
            arith_in_col_17_d5 <=  arith_in_col_17_d4;
            arith_in_col_17_d6 <=  arith_in_col_17_d5;
            arith_in_col_17_d7 <=  arith_in_col_17_d6;
            arith_in_col_17_d8 <=  arith_in_col_17_d7;
            arith_in_col_17_d9 <=  arith_in_col_17_d8;
            arith_in_col_17_d10 <=  arith_in_col_17_d9;
            arith_in_col_17_d11 <=  arith_in_col_17_d10;
            arith_in_col_17_d12 <=  arith_in_col_17_d11;
            arith_in_col_17_d13 <=  arith_in_col_17_d12;
            arith_in_col_17_d14 <=  arith_in_col_17_d13;
            arith_in_col_17_d15 <=  arith_in_col_17_d14;
            arith_in_col_17_d16 <=  arith_in_col_17_d15;
            arith_in_col_17_d17 <=  arith_in_col_17_d16;
            arith_in_col_18_d1 <=  arith_in_col_18;
            arith_in_col_18_d2 <=  arith_in_col_18_d1;
            arith_in_col_18_d3 <=  arith_in_col_18_d2;
            arith_in_col_18_d4 <=  arith_in_col_18_d3;
            arith_in_col_18_d5 <=  arith_in_col_18_d4;
            arith_in_col_18_d6 <=  arith_in_col_18_d5;
            arith_in_col_18_d7 <=  arith_in_col_18_d6;
            arith_in_col_18_d8 <=  arith_in_col_18_d7;
            arith_in_col_18_d9 <=  arith_in_col_18_d8;
            arith_in_col_18_d10 <=  arith_in_col_18_d9;
            arith_in_col_18_d11 <=  arith_in_col_18_d10;
            arith_in_col_18_d12 <=  arith_in_col_18_d11;
            arith_in_col_18_d13 <=  arith_in_col_18_d12;
            arith_in_col_18_d14 <=  arith_in_col_18_d13;
            arith_in_col_18_d15 <=  arith_in_col_18_d14;
            arith_in_col_18_d16 <=  arith_in_col_18_d15;
            arith_in_col_18_d17 <=  arith_in_col_18_d16;
            arith_in_col_18_d18 <=  arith_in_col_18_d17;
            arith_in_col_19_d1 <=  arith_in_col_19;
            arith_in_col_19_d2 <=  arith_in_col_19_d1;
            arith_in_col_19_d3 <=  arith_in_col_19_d2;
            arith_in_col_19_d4 <=  arith_in_col_19_d3;
            arith_in_col_19_d5 <=  arith_in_col_19_d4;
            arith_in_col_19_d6 <=  arith_in_col_19_d5;
            arith_in_col_19_d7 <=  arith_in_col_19_d6;
            arith_in_col_19_d8 <=  arith_in_col_19_d7;
            arith_in_col_19_d9 <=  arith_in_col_19_d8;
            arith_in_col_19_d10 <=  arith_in_col_19_d9;
            arith_in_col_19_d11 <=  arith_in_col_19_d10;
            arith_in_col_19_d12 <=  arith_in_col_19_d11;
            arith_in_col_19_d13 <=  arith_in_col_19_d12;
            arith_in_col_19_d14 <=  arith_in_col_19_d13;
            arith_in_col_19_d15 <=  arith_in_col_19_d14;
            arith_in_col_19_d16 <=  arith_in_col_19_d15;
            arith_in_col_19_d17 <=  arith_in_col_19_d16;
            arith_in_col_19_d18 <=  arith_in_col_19_d17;
            arith_in_col_19_d19 <=  arith_in_col_19_d18;
            arith_in_col_20_d1 <=  arith_in_col_20;
            arith_in_col_20_d2 <=  arith_in_col_20_d1;
            arith_in_col_20_d3 <=  arith_in_col_20_d2;
            arith_in_col_20_d4 <=  arith_in_col_20_d3;
            arith_in_col_20_d5 <=  arith_in_col_20_d4;
            arith_in_col_20_d6 <=  arith_in_col_20_d5;
            arith_in_col_20_d7 <=  arith_in_col_20_d6;
            arith_in_col_20_d8 <=  arith_in_col_20_d7;
            arith_in_col_20_d9 <=  arith_in_col_20_d8;
            arith_in_col_20_d10 <=  arith_in_col_20_d9;
            arith_in_col_20_d11 <=  arith_in_col_20_d10;
            arith_in_col_20_d12 <=  arith_in_col_20_d11;
            arith_in_col_20_d13 <=  arith_in_col_20_d12;
            arith_in_col_20_d14 <=  arith_in_col_20_d13;
            arith_in_col_20_d15 <=  arith_in_col_20_d14;
            arith_in_col_20_d16 <=  arith_in_col_20_d15;
            arith_in_col_20_d17 <=  arith_in_col_20_d16;
            arith_in_col_20_d18 <=  arith_in_col_20_d17;
            arith_in_col_20_d19 <=  arith_in_col_20_d18;
            arith_in_col_20_d20 <=  arith_in_col_20_d19;
            arith_in_col_21_d1 <=  arith_in_col_21;
            arith_in_col_21_d2 <=  arith_in_col_21_d1;
            arith_in_col_21_d3 <=  arith_in_col_21_d2;
            arith_in_col_21_d4 <=  arith_in_col_21_d3;
            arith_in_col_21_d5 <=  arith_in_col_21_d4;
            arith_in_col_21_d6 <=  arith_in_col_21_d5;
            arith_in_col_21_d7 <=  arith_in_col_21_d6;
            arith_in_col_21_d8 <=  arith_in_col_21_d7;
            arith_in_col_21_d9 <=  arith_in_col_21_d8;
            arith_in_col_21_d10 <=  arith_in_col_21_d9;
            arith_in_col_21_d11 <=  arith_in_col_21_d10;
            arith_in_col_21_d12 <=  arith_in_col_21_d11;
            arith_in_col_21_d13 <=  arith_in_col_21_d12;
            arith_in_col_21_d14 <=  arith_in_col_21_d13;
            arith_in_col_21_d15 <=  arith_in_col_21_d14;
            arith_in_col_21_d16 <=  arith_in_col_21_d15;
            arith_in_col_21_d17 <=  arith_in_col_21_d16;
            arith_in_col_21_d18 <=  arith_in_col_21_d17;
            arith_in_col_21_d19 <=  arith_in_col_21_d18;
            arith_in_col_21_d20 <=  arith_in_col_21_d19;
            arith_in_col_21_d21 <=  arith_in_col_21_d20;
            arith_in_col_22_d1 <=  arith_in_col_22;
            arith_in_col_22_d2 <=  arith_in_col_22_d1;
            arith_in_col_22_d3 <=  arith_in_col_22_d2;
            arith_in_col_22_d4 <=  arith_in_col_22_d3;
            arith_in_col_22_d5 <=  arith_in_col_22_d4;
            arith_in_col_22_d6 <=  arith_in_col_22_d5;
            arith_in_col_22_d7 <=  arith_in_col_22_d6;
            arith_in_col_22_d8 <=  arith_in_col_22_d7;
            arith_in_col_22_d9 <=  arith_in_col_22_d8;
            arith_in_col_22_d10 <=  arith_in_col_22_d9;
            arith_in_col_22_d11 <=  arith_in_col_22_d10;
            arith_in_col_22_d12 <=  arith_in_col_22_d11;
            arith_in_col_22_d13 <=  arith_in_col_22_d12;
            arith_in_col_22_d14 <=  arith_in_col_22_d13;
            arith_in_col_22_d15 <=  arith_in_col_22_d14;
            arith_in_col_22_d16 <=  arith_in_col_22_d15;
            arith_in_col_22_d17 <=  arith_in_col_22_d16;
            arith_in_col_22_d18 <=  arith_in_col_22_d17;
            arith_in_col_22_d19 <=  arith_in_col_22_d18;
            arith_in_col_22_d20 <=  arith_in_col_22_d19;
            arith_in_col_22_d21 <=  arith_in_col_22_d20;
            arith_in_col_22_d22 <=  arith_in_col_22_d21;
            arith_in_col_23_d1 <=  arith_in_col_23;
            arith_in_col_23_d2 <=  arith_in_col_23_d1;
            arith_in_col_23_d3 <=  arith_in_col_23_d2;
            arith_in_col_23_d4 <=  arith_in_col_23_d3;
            arith_in_col_23_d5 <=  arith_in_col_23_d4;
            arith_in_col_23_d6 <=  arith_in_col_23_d5;
            arith_in_col_23_d7 <=  arith_in_col_23_d6;
            arith_in_col_23_d8 <=  arith_in_col_23_d7;
            arith_in_col_23_d9 <=  arith_in_col_23_d8;
            arith_in_col_23_d10 <=  arith_in_col_23_d9;
            arith_in_col_23_d11 <=  arith_in_col_23_d10;
            arith_in_col_23_d12 <=  arith_in_col_23_d11;
            arith_in_col_23_d13 <=  arith_in_col_23_d12;
            arith_in_col_23_d14 <=  arith_in_col_23_d13;
            arith_in_col_23_d15 <=  arith_in_col_23_d14;
            arith_in_col_23_d16 <=  arith_in_col_23_d15;
            arith_in_col_23_d17 <=  arith_in_col_23_d16;
            arith_in_col_23_d18 <=  arith_in_col_23_d17;
            arith_in_col_23_d19 <=  arith_in_col_23_d18;
            arith_in_col_23_d20 <=  arith_in_col_23_d19;
            arith_in_col_23_d21 <=  arith_in_col_23_d20;
            arith_in_col_23_d22 <=  arith_in_col_23_d21;
            arith_in_col_23_d23 <=  arith_in_col_23_d22;
            arith_in_col_24_d1 <=  arith_in_col_24;
            arith_in_col_24_d2 <=  arith_in_col_24_d1;
            arith_in_col_24_d3 <=  arith_in_col_24_d2;
            arith_in_col_24_d4 <=  arith_in_col_24_d3;
            arith_in_col_24_d5 <=  arith_in_col_24_d4;
            arith_in_col_24_d6 <=  arith_in_col_24_d5;
            arith_in_col_24_d7 <=  arith_in_col_24_d6;
            arith_in_col_24_d8 <=  arith_in_col_24_d7;
            arith_in_col_24_d9 <=  arith_in_col_24_d8;
            arith_in_col_24_d10 <=  arith_in_col_24_d9;
            arith_in_col_24_d11 <=  arith_in_col_24_d10;
            arith_in_col_24_d12 <=  arith_in_col_24_d11;
            arith_in_col_24_d13 <=  arith_in_col_24_d12;
            arith_in_col_24_d14 <=  arith_in_col_24_d13;
            arith_in_col_24_d15 <=  arith_in_col_24_d14;
            arith_in_col_24_d16 <=  arith_in_col_24_d15;
            arith_in_col_24_d17 <=  arith_in_col_24_d16;
            arith_in_col_24_d18 <=  arith_in_col_24_d17;
            arith_in_col_24_d19 <=  arith_in_col_24_d18;
            arith_in_col_24_d20 <=  arith_in_col_24_d19;
            arith_in_col_24_d21 <=  arith_in_col_24_d20;
            arith_in_col_24_d22 <=  arith_in_col_24_d21;
            arith_in_col_24_d23 <=  arith_in_col_24_d22;
            arith_in_col_24_d24 <=  arith_in_col_24_d23;
            arith_in_col_25_d1 <=  arith_in_col_25;
            arith_in_col_25_d2 <=  arith_in_col_25_d1;
            arith_in_col_25_d3 <=  arith_in_col_25_d2;
            arith_in_col_25_d4 <=  arith_in_col_25_d3;
            arith_in_col_25_d5 <=  arith_in_col_25_d4;
            arith_in_col_25_d6 <=  arith_in_col_25_d5;
            arith_in_col_25_d7 <=  arith_in_col_25_d6;
            arith_in_col_25_d8 <=  arith_in_col_25_d7;
            arith_in_col_25_d9 <=  arith_in_col_25_d8;
            arith_in_col_25_d10 <=  arith_in_col_25_d9;
            arith_in_col_25_d11 <=  arith_in_col_25_d10;
            arith_in_col_25_d12 <=  arith_in_col_25_d11;
            arith_in_col_25_d13 <=  arith_in_col_25_d12;
            arith_in_col_25_d14 <=  arith_in_col_25_d13;
            arith_in_col_25_d15 <=  arith_in_col_25_d14;
            arith_in_col_25_d16 <=  arith_in_col_25_d15;
            arith_in_col_25_d17 <=  arith_in_col_25_d16;
            arith_in_col_25_d18 <=  arith_in_col_25_d17;
            arith_in_col_25_d19 <=  arith_in_col_25_d18;
            arith_in_col_25_d20 <=  arith_in_col_25_d19;
            arith_in_col_25_d21 <=  arith_in_col_25_d20;
            arith_in_col_25_d22 <=  arith_in_col_25_d21;
            arith_in_col_25_d23 <=  arith_in_col_25_d22;
            arith_in_col_25_d24 <=  arith_in_col_25_d23;
            arith_in_col_25_d25 <=  arith_in_col_25_d24;
            arith_in_col_26_d1 <=  arith_in_col_26;
            arith_in_col_26_d2 <=  arith_in_col_26_d1;
            arith_in_col_26_d3 <=  arith_in_col_26_d2;
            arith_in_col_26_d4 <=  arith_in_col_26_d3;
            arith_in_col_26_d5 <=  arith_in_col_26_d4;
            arith_in_col_26_d6 <=  arith_in_col_26_d5;
            arith_in_col_26_d7 <=  arith_in_col_26_d6;
            arith_in_col_26_d8 <=  arith_in_col_26_d7;
            arith_in_col_26_d9 <=  arith_in_col_26_d8;
            arith_in_col_26_d10 <=  arith_in_col_26_d9;
            arith_in_col_26_d11 <=  arith_in_col_26_d10;
            arith_in_col_26_d12 <=  arith_in_col_26_d11;
            arith_in_col_26_d13 <=  arith_in_col_26_d12;
            arith_in_col_26_d14 <=  arith_in_col_26_d13;
            arith_in_col_26_d15 <=  arith_in_col_26_d14;
            arith_in_col_26_d16 <=  arith_in_col_26_d15;
            arith_in_col_26_d17 <=  arith_in_col_26_d16;
            arith_in_col_26_d18 <=  arith_in_col_26_d17;
            arith_in_col_26_d19 <=  arith_in_col_26_d18;
            arith_in_col_26_d20 <=  arith_in_col_26_d19;
            arith_in_col_26_d21 <=  arith_in_col_26_d20;
            arith_in_col_26_d22 <=  arith_in_col_26_d21;
            arith_in_col_26_d23 <=  arith_in_col_26_d22;
            arith_in_col_26_d24 <=  arith_in_col_26_d23;
            arith_in_col_26_d25 <=  arith_in_col_26_d24;
            arith_in_col_26_d26 <=  arith_in_col_26_d25;
            arith_in_col_27_d1 <=  arith_in_col_27;
            arith_in_col_27_d2 <=  arith_in_col_27_d1;
            arith_in_col_27_d3 <=  arith_in_col_27_d2;
            arith_in_col_27_d4 <=  arith_in_col_27_d3;
            arith_in_col_27_d5 <=  arith_in_col_27_d4;
            arith_in_col_27_d6 <=  arith_in_col_27_d5;
            arith_in_col_27_d7 <=  arith_in_col_27_d6;
            arith_in_col_27_d8 <=  arith_in_col_27_d7;
            arith_in_col_27_d9 <=  arith_in_col_27_d8;
            arith_in_col_27_d10 <=  arith_in_col_27_d9;
            arith_in_col_27_d11 <=  arith_in_col_27_d10;
            arith_in_col_27_d12 <=  arith_in_col_27_d11;
            arith_in_col_27_d13 <=  arith_in_col_27_d12;
            arith_in_col_27_d14 <=  arith_in_col_27_d13;
            arith_in_col_27_d15 <=  arith_in_col_27_d14;
            arith_in_col_27_d16 <=  arith_in_col_27_d15;
            arith_in_col_27_d17 <=  arith_in_col_27_d16;
            arith_in_col_27_d18 <=  arith_in_col_27_d17;
            arith_in_col_27_d19 <=  arith_in_col_27_d18;
            arith_in_col_27_d20 <=  arith_in_col_27_d19;
            arith_in_col_27_d21 <=  arith_in_col_27_d20;
            arith_in_col_27_d22 <=  arith_in_col_27_d21;
            arith_in_col_27_d23 <=  arith_in_col_27_d22;
            arith_in_col_27_d24 <=  arith_in_col_27_d23;
            arith_in_col_27_d25 <=  arith_in_col_27_d24;
            arith_in_col_27_d26 <=  arith_in_col_27_d25;
            arith_in_col_27_d27 <=  arith_in_col_27_d26;
            arith_in_col_28_d1 <=  arith_in_col_28;
            arith_in_col_28_d2 <=  arith_in_col_28_d1;
            arith_in_col_28_d3 <=  arith_in_col_28_d2;
            arith_in_col_28_d4 <=  arith_in_col_28_d3;
            arith_in_col_28_d5 <=  arith_in_col_28_d4;
            arith_in_col_28_d6 <=  arith_in_col_28_d5;
            arith_in_col_28_d7 <=  arith_in_col_28_d6;
            arith_in_col_28_d8 <=  arith_in_col_28_d7;
            arith_in_col_28_d9 <=  arith_in_col_28_d8;
            arith_in_col_28_d10 <=  arith_in_col_28_d9;
            arith_in_col_28_d11 <=  arith_in_col_28_d10;
            arith_in_col_28_d12 <=  arith_in_col_28_d11;
            arith_in_col_28_d13 <=  arith_in_col_28_d12;
            arith_in_col_28_d14 <=  arith_in_col_28_d13;
            arith_in_col_28_d15 <=  arith_in_col_28_d14;
            arith_in_col_28_d16 <=  arith_in_col_28_d15;
            arith_in_col_28_d17 <=  arith_in_col_28_d16;
            arith_in_col_28_d18 <=  arith_in_col_28_d17;
            arith_in_col_28_d19 <=  arith_in_col_28_d18;
            arith_in_col_28_d20 <=  arith_in_col_28_d19;
            arith_in_col_28_d21 <=  arith_in_col_28_d20;
            arith_in_col_28_d22 <=  arith_in_col_28_d21;
            arith_in_col_28_d23 <=  arith_in_col_28_d22;
            arith_in_col_28_d24 <=  arith_in_col_28_d23;
            arith_in_col_28_d25 <=  arith_in_col_28_d24;
            arith_in_col_28_d26 <=  arith_in_col_28_d25;
            arith_in_col_28_d27 <=  arith_in_col_28_d26;
            arith_in_col_28_d28 <=  arith_in_col_28_d27;
            arith_in_col_29_d1 <=  arith_in_col_29;
            arith_in_col_29_d2 <=  arith_in_col_29_d1;
            arith_in_col_29_d3 <=  arith_in_col_29_d2;
            arith_in_col_29_d4 <=  arith_in_col_29_d3;
            arith_in_col_29_d5 <=  arith_in_col_29_d4;
            arith_in_col_29_d6 <=  arith_in_col_29_d5;
            arith_in_col_29_d7 <=  arith_in_col_29_d6;
            arith_in_col_29_d8 <=  arith_in_col_29_d7;
            arith_in_col_29_d9 <=  arith_in_col_29_d8;
            arith_in_col_29_d10 <=  arith_in_col_29_d9;
            arith_in_col_29_d11 <=  arith_in_col_29_d10;
            arith_in_col_29_d12 <=  arith_in_col_29_d11;
            arith_in_col_29_d13 <=  arith_in_col_29_d12;
            arith_in_col_29_d14 <=  arith_in_col_29_d13;
            arith_in_col_29_d15 <=  arith_in_col_29_d14;
            arith_in_col_29_d16 <=  arith_in_col_29_d15;
            arith_in_col_29_d17 <=  arith_in_col_29_d16;
            arith_in_col_29_d18 <=  arith_in_col_29_d17;
            arith_in_col_29_d19 <=  arith_in_col_29_d18;
            arith_in_col_29_d20 <=  arith_in_col_29_d19;
            arith_in_col_29_d21 <=  arith_in_col_29_d20;
            arith_in_col_29_d22 <=  arith_in_col_29_d21;
            arith_in_col_29_d23 <=  arith_in_col_29_d22;
            arith_in_col_29_d24 <=  arith_in_col_29_d23;
            arith_in_col_29_d25 <=  arith_in_col_29_d24;
            arith_in_col_29_d26 <=  arith_in_col_29_d25;
            arith_in_col_29_d27 <=  arith_in_col_29_d26;
            arith_in_col_29_d28 <=  arith_in_col_29_d27;
            arith_in_col_29_d29 <=  arith_in_col_29_d28;
            arith_in_col_30_d1 <=  arith_in_col_30;
            arith_in_col_30_d2 <=  arith_in_col_30_d1;
            arith_in_col_30_d3 <=  arith_in_col_30_d2;
            arith_in_col_30_d4 <=  arith_in_col_30_d3;
            arith_in_col_30_d5 <=  arith_in_col_30_d4;
            arith_in_col_30_d6 <=  arith_in_col_30_d5;
            arith_in_col_30_d7 <=  arith_in_col_30_d6;
            arith_in_col_30_d8 <=  arith_in_col_30_d7;
            arith_in_col_30_d9 <=  arith_in_col_30_d8;
            arith_in_col_30_d10 <=  arith_in_col_30_d9;
            arith_in_col_30_d11 <=  arith_in_col_30_d10;
            arith_in_col_30_d12 <=  arith_in_col_30_d11;
            arith_in_col_30_d13 <=  arith_in_col_30_d12;
            arith_in_col_30_d14 <=  arith_in_col_30_d13;
            arith_in_col_30_d15 <=  arith_in_col_30_d14;
            arith_in_col_30_d16 <=  arith_in_col_30_d15;
            arith_in_col_30_d17 <=  arith_in_col_30_d16;
            arith_in_col_30_d18 <=  arith_in_col_30_d17;
            arith_in_col_30_d19 <=  arith_in_col_30_d18;
            arith_in_col_30_d20 <=  arith_in_col_30_d19;
            arith_in_col_30_d21 <=  arith_in_col_30_d20;
            arith_in_col_30_d22 <=  arith_in_col_30_d21;
            arith_in_col_30_d23 <=  arith_in_col_30_d22;
            arith_in_col_30_d24 <=  arith_in_col_30_d23;
            arith_in_col_30_d25 <=  arith_in_col_30_d24;
            arith_in_col_30_d26 <=  arith_in_col_30_d25;
            arith_in_col_30_d27 <=  arith_in_col_30_d26;
            arith_in_col_30_d28 <=  arith_in_col_30_d27;
            arith_in_col_30_d29 <=  arith_in_col_30_d28;
            arith_in_col_30_d30 <=  arith_in_col_30_d29;
            arith_out_col_out_0_d1 <=  arith_out_col_out_0;
            arith_out_col_out_0_d2 <=  arith_out_col_out_0_d1;
            arith_out_col_out_0_d3 <=  arith_out_col_out_0_d2;
            arith_out_col_out_0_d4 <=  arith_out_col_out_0_d3;
            arith_out_col_out_0_d5 <=  arith_out_col_out_0_d4;
            arith_out_col_out_0_d6 <=  arith_out_col_out_0_d5;
            arith_out_col_out_0_d7 <=  arith_out_col_out_0_d6;
            arith_out_col_out_0_d8 <=  arith_out_col_out_0_d7;
            arith_out_col_out_0_d9 <=  arith_out_col_out_0_d8;
            arith_out_col_out_0_d10 <=  arith_out_col_out_0_d9;
            arith_out_col_out_0_d11 <=  arith_out_col_out_0_d10;
            arith_out_col_out_0_d12 <=  arith_out_col_out_0_d11;
            arith_out_col_out_0_d13 <=  arith_out_col_out_0_d12;
            arith_out_col_out_0_d14 <=  arith_out_col_out_0_d13;
            arith_out_col_out_0_d15 <=  arith_out_col_out_0_d14;
            arith_out_col_out_0_d16 <=  arith_out_col_out_0_d15;
            arith_out_col_out_0_d17 <=  arith_out_col_out_0_d16;
            arith_out_col_out_0_d18 <=  arith_out_col_out_0_d17;
            arith_out_col_out_0_d19 <=  arith_out_col_out_0_d18;
            arith_out_col_out_0_d20 <=  arith_out_col_out_0_d19;
            arith_out_col_out_0_d21 <=  arith_out_col_out_0_d20;
            arith_out_col_out_0_d22 <=  arith_out_col_out_0_d21;
            arith_out_col_out_0_d23 <=  arith_out_col_out_0_d22;
            arith_out_col_out_0_d24 <=  arith_out_col_out_0_d23;
            arith_out_col_out_0_d25 <=  arith_out_col_out_0_d24;
            arith_out_col_out_0_d26 <=  arith_out_col_out_0_d25;
            arith_out_col_out_0_d27 <=  arith_out_col_out_0_d26;
            arith_out_col_out_0_d28 <=  arith_out_col_out_0_d27;
            arith_out_col_out_0_d29 <=  arith_out_col_out_0_d28;
            arith_out_col_out_0_d30 <=  arith_out_col_out_0_d29;
            arith_out_col_out_1_d1 <=  arith_out_col_out_1;
            arith_out_col_out_1_d2 <=  arith_out_col_out_1_d1;
            arith_out_col_out_1_d3 <=  arith_out_col_out_1_d2;
            arith_out_col_out_1_d4 <=  arith_out_col_out_1_d3;
            arith_out_col_out_1_d5 <=  arith_out_col_out_1_d4;
            arith_out_col_out_1_d6 <=  arith_out_col_out_1_d5;
            arith_out_col_out_1_d7 <=  arith_out_col_out_1_d6;
            arith_out_col_out_1_d8 <=  arith_out_col_out_1_d7;
            arith_out_col_out_1_d9 <=  arith_out_col_out_1_d8;
            arith_out_col_out_1_d10 <=  arith_out_col_out_1_d9;
            arith_out_col_out_1_d11 <=  arith_out_col_out_1_d10;
            arith_out_col_out_1_d12 <=  arith_out_col_out_1_d11;
            arith_out_col_out_1_d13 <=  arith_out_col_out_1_d12;
            arith_out_col_out_1_d14 <=  arith_out_col_out_1_d13;
            arith_out_col_out_1_d15 <=  arith_out_col_out_1_d14;
            arith_out_col_out_1_d16 <=  arith_out_col_out_1_d15;
            arith_out_col_out_1_d17 <=  arith_out_col_out_1_d16;
            arith_out_col_out_1_d18 <=  arith_out_col_out_1_d17;
            arith_out_col_out_1_d19 <=  arith_out_col_out_1_d18;
            arith_out_col_out_1_d20 <=  arith_out_col_out_1_d19;
            arith_out_col_out_1_d21 <=  arith_out_col_out_1_d20;
            arith_out_col_out_1_d22 <=  arith_out_col_out_1_d21;
            arith_out_col_out_1_d23 <=  arith_out_col_out_1_d22;
            arith_out_col_out_1_d24 <=  arith_out_col_out_1_d23;
            arith_out_col_out_1_d25 <=  arith_out_col_out_1_d24;
            arith_out_col_out_1_d26 <=  arith_out_col_out_1_d25;
            arith_out_col_out_1_d27 <=  arith_out_col_out_1_d26;
            arith_out_col_out_1_d28 <=  arith_out_col_out_1_d27;
            arith_out_col_out_1_d29 <=  arith_out_col_out_1_d28;
            arith_out_col_out_2_d1 <=  arith_out_col_out_2;
            arith_out_col_out_2_d2 <=  arith_out_col_out_2_d1;
            arith_out_col_out_2_d3 <=  arith_out_col_out_2_d2;
            arith_out_col_out_2_d4 <=  arith_out_col_out_2_d3;
            arith_out_col_out_2_d5 <=  arith_out_col_out_2_d4;
            arith_out_col_out_2_d6 <=  arith_out_col_out_2_d5;
            arith_out_col_out_2_d7 <=  arith_out_col_out_2_d6;
            arith_out_col_out_2_d8 <=  arith_out_col_out_2_d7;
            arith_out_col_out_2_d9 <=  arith_out_col_out_2_d8;
            arith_out_col_out_2_d10 <=  arith_out_col_out_2_d9;
            arith_out_col_out_2_d11 <=  arith_out_col_out_2_d10;
            arith_out_col_out_2_d12 <=  arith_out_col_out_2_d11;
            arith_out_col_out_2_d13 <=  arith_out_col_out_2_d12;
            arith_out_col_out_2_d14 <=  arith_out_col_out_2_d13;
            arith_out_col_out_2_d15 <=  arith_out_col_out_2_d14;
            arith_out_col_out_2_d16 <=  arith_out_col_out_2_d15;
            arith_out_col_out_2_d17 <=  arith_out_col_out_2_d16;
            arith_out_col_out_2_d18 <=  arith_out_col_out_2_d17;
            arith_out_col_out_2_d19 <=  arith_out_col_out_2_d18;
            arith_out_col_out_2_d20 <=  arith_out_col_out_2_d19;
            arith_out_col_out_2_d21 <=  arith_out_col_out_2_d20;
            arith_out_col_out_2_d22 <=  arith_out_col_out_2_d21;
            arith_out_col_out_2_d23 <=  arith_out_col_out_2_d22;
            arith_out_col_out_2_d24 <=  arith_out_col_out_2_d23;
            arith_out_col_out_2_d25 <=  arith_out_col_out_2_d24;
            arith_out_col_out_2_d26 <=  arith_out_col_out_2_d25;
            arith_out_col_out_2_d27 <=  arith_out_col_out_2_d26;
            arith_out_col_out_2_d28 <=  arith_out_col_out_2_d27;
            arith_out_col_out_3_d1 <=  arith_out_col_out_3;
            arith_out_col_out_3_d2 <=  arith_out_col_out_3_d1;
            arith_out_col_out_3_d3 <=  arith_out_col_out_3_d2;
            arith_out_col_out_3_d4 <=  arith_out_col_out_3_d3;
            arith_out_col_out_3_d5 <=  arith_out_col_out_3_d4;
            arith_out_col_out_3_d6 <=  arith_out_col_out_3_d5;
            arith_out_col_out_3_d7 <=  arith_out_col_out_3_d6;
            arith_out_col_out_3_d8 <=  arith_out_col_out_3_d7;
            arith_out_col_out_3_d9 <=  arith_out_col_out_3_d8;
            arith_out_col_out_3_d10 <=  arith_out_col_out_3_d9;
            arith_out_col_out_3_d11 <=  arith_out_col_out_3_d10;
            arith_out_col_out_3_d12 <=  arith_out_col_out_3_d11;
            arith_out_col_out_3_d13 <=  arith_out_col_out_3_d12;
            arith_out_col_out_3_d14 <=  arith_out_col_out_3_d13;
            arith_out_col_out_3_d15 <=  arith_out_col_out_3_d14;
            arith_out_col_out_3_d16 <=  arith_out_col_out_3_d15;
            arith_out_col_out_3_d17 <=  arith_out_col_out_3_d16;
            arith_out_col_out_3_d18 <=  arith_out_col_out_3_d17;
            arith_out_col_out_3_d19 <=  arith_out_col_out_3_d18;
            arith_out_col_out_3_d20 <=  arith_out_col_out_3_d19;
            arith_out_col_out_3_d21 <=  arith_out_col_out_3_d20;
            arith_out_col_out_3_d22 <=  arith_out_col_out_3_d21;
            arith_out_col_out_3_d23 <=  arith_out_col_out_3_d22;
            arith_out_col_out_3_d24 <=  arith_out_col_out_3_d23;
            arith_out_col_out_3_d25 <=  arith_out_col_out_3_d24;
            arith_out_col_out_3_d26 <=  arith_out_col_out_3_d25;
            arith_out_col_out_3_d27 <=  arith_out_col_out_3_d26;
            arith_out_col_out_4_d1 <=  arith_out_col_out_4;
            arith_out_col_out_4_d2 <=  arith_out_col_out_4_d1;
            arith_out_col_out_4_d3 <=  arith_out_col_out_4_d2;
            arith_out_col_out_4_d4 <=  arith_out_col_out_4_d3;
            arith_out_col_out_4_d5 <=  arith_out_col_out_4_d4;
            arith_out_col_out_4_d6 <=  arith_out_col_out_4_d5;
            arith_out_col_out_4_d7 <=  arith_out_col_out_4_d6;
            arith_out_col_out_4_d8 <=  arith_out_col_out_4_d7;
            arith_out_col_out_4_d9 <=  arith_out_col_out_4_d8;
            arith_out_col_out_4_d10 <=  arith_out_col_out_4_d9;
            arith_out_col_out_4_d11 <=  arith_out_col_out_4_d10;
            arith_out_col_out_4_d12 <=  arith_out_col_out_4_d11;
            arith_out_col_out_4_d13 <=  arith_out_col_out_4_d12;
            arith_out_col_out_4_d14 <=  arith_out_col_out_4_d13;
            arith_out_col_out_4_d15 <=  arith_out_col_out_4_d14;
            arith_out_col_out_4_d16 <=  arith_out_col_out_4_d15;
            arith_out_col_out_4_d17 <=  arith_out_col_out_4_d16;
            arith_out_col_out_4_d18 <=  arith_out_col_out_4_d17;
            arith_out_col_out_4_d19 <=  arith_out_col_out_4_d18;
            arith_out_col_out_4_d20 <=  arith_out_col_out_4_d19;
            arith_out_col_out_4_d21 <=  arith_out_col_out_4_d20;
            arith_out_col_out_4_d22 <=  arith_out_col_out_4_d21;
            arith_out_col_out_4_d23 <=  arith_out_col_out_4_d22;
            arith_out_col_out_4_d24 <=  arith_out_col_out_4_d23;
            arith_out_col_out_4_d25 <=  arith_out_col_out_4_d24;
            arith_out_col_out_4_d26 <=  arith_out_col_out_4_d25;
            arith_out_col_out_5_d1 <=  arith_out_col_out_5;
            arith_out_col_out_5_d2 <=  arith_out_col_out_5_d1;
            arith_out_col_out_5_d3 <=  arith_out_col_out_5_d2;
            arith_out_col_out_5_d4 <=  arith_out_col_out_5_d3;
            arith_out_col_out_5_d5 <=  arith_out_col_out_5_d4;
            arith_out_col_out_5_d6 <=  arith_out_col_out_5_d5;
            arith_out_col_out_5_d7 <=  arith_out_col_out_5_d6;
            arith_out_col_out_5_d8 <=  arith_out_col_out_5_d7;
            arith_out_col_out_5_d9 <=  arith_out_col_out_5_d8;
            arith_out_col_out_5_d10 <=  arith_out_col_out_5_d9;
            arith_out_col_out_5_d11 <=  arith_out_col_out_5_d10;
            arith_out_col_out_5_d12 <=  arith_out_col_out_5_d11;
            arith_out_col_out_5_d13 <=  arith_out_col_out_5_d12;
            arith_out_col_out_5_d14 <=  arith_out_col_out_5_d13;
            arith_out_col_out_5_d15 <=  arith_out_col_out_5_d14;
            arith_out_col_out_5_d16 <=  arith_out_col_out_5_d15;
            arith_out_col_out_5_d17 <=  arith_out_col_out_5_d16;
            arith_out_col_out_5_d18 <=  arith_out_col_out_5_d17;
            arith_out_col_out_5_d19 <=  arith_out_col_out_5_d18;
            arith_out_col_out_5_d20 <=  arith_out_col_out_5_d19;
            arith_out_col_out_5_d21 <=  arith_out_col_out_5_d20;
            arith_out_col_out_5_d22 <=  arith_out_col_out_5_d21;
            arith_out_col_out_5_d23 <=  arith_out_col_out_5_d22;
            arith_out_col_out_5_d24 <=  arith_out_col_out_5_d23;
            arith_out_col_out_5_d25 <=  arith_out_col_out_5_d24;
            arith_out_col_out_6_d1 <=  arith_out_col_out_6;
            arith_out_col_out_6_d2 <=  arith_out_col_out_6_d1;
            arith_out_col_out_6_d3 <=  arith_out_col_out_6_d2;
            arith_out_col_out_6_d4 <=  arith_out_col_out_6_d3;
            arith_out_col_out_6_d5 <=  arith_out_col_out_6_d4;
            arith_out_col_out_6_d6 <=  arith_out_col_out_6_d5;
            arith_out_col_out_6_d7 <=  arith_out_col_out_6_d6;
            arith_out_col_out_6_d8 <=  arith_out_col_out_6_d7;
            arith_out_col_out_6_d9 <=  arith_out_col_out_6_d8;
            arith_out_col_out_6_d10 <=  arith_out_col_out_6_d9;
            arith_out_col_out_6_d11 <=  arith_out_col_out_6_d10;
            arith_out_col_out_6_d12 <=  arith_out_col_out_6_d11;
            arith_out_col_out_6_d13 <=  arith_out_col_out_6_d12;
            arith_out_col_out_6_d14 <=  arith_out_col_out_6_d13;
            arith_out_col_out_6_d15 <=  arith_out_col_out_6_d14;
            arith_out_col_out_6_d16 <=  arith_out_col_out_6_d15;
            arith_out_col_out_6_d17 <=  arith_out_col_out_6_d16;
            arith_out_col_out_6_d18 <=  arith_out_col_out_6_d17;
            arith_out_col_out_6_d19 <=  arith_out_col_out_6_d18;
            arith_out_col_out_6_d20 <=  arith_out_col_out_6_d19;
            arith_out_col_out_6_d21 <=  arith_out_col_out_6_d20;
            arith_out_col_out_6_d22 <=  arith_out_col_out_6_d21;
            arith_out_col_out_6_d23 <=  arith_out_col_out_6_d22;
            arith_out_col_out_6_d24 <=  arith_out_col_out_6_d23;
            arith_out_col_out_7_d1 <=  arith_out_col_out_7;
            arith_out_col_out_7_d2 <=  arith_out_col_out_7_d1;
            arith_out_col_out_7_d3 <=  arith_out_col_out_7_d2;
            arith_out_col_out_7_d4 <=  arith_out_col_out_7_d3;
            arith_out_col_out_7_d5 <=  arith_out_col_out_7_d4;
            arith_out_col_out_7_d6 <=  arith_out_col_out_7_d5;
            arith_out_col_out_7_d7 <=  arith_out_col_out_7_d6;
            arith_out_col_out_7_d8 <=  arith_out_col_out_7_d7;
            arith_out_col_out_7_d9 <=  arith_out_col_out_7_d8;
            arith_out_col_out_7_d10 <=  arith_out_col_out_7_d9;
            arith_out_col_out_7_d11 <=  arith_out_col_out_7_d10;
            arith_out_col_out_7_d12 <=  arith_out_col_out_7_d11;
            arith_out_col_out_7_d13 <=  arith_out_col_out_7_d12;
            arith_out_col_out_7_d14 <=  arith_out_col_out_7_d13;
            arith_out_col_out_7_d15 <=  arith_out_col_out_7_d14;
            arith_out_col_out_7_d16 <=  arith_out_col_out_7_d15;
            arith_out_col_out_7_d17 <=  arith_out_col_out_7_d16;
            arith_out_col_out_7_d18 <=  arith_out_col_out_7_d17;
            arith_out_col_out_7_d19 <=  arith_out_col_out_7_d18;
            arith_out_col_out_7_d20 <=  arith_out_col_out_7_d19;
            arith_out_col_out_7_d21 <=  arith_out_col_out_7_d20;
            arith_out_col_out_7_d22 <=  arith_out_col_out_7_d21;
            arith_out_col_out_7_d23 <=  arith_out_col_out_7_d22;
            arith_out_col_out_8_d1 <=  arith_out_col_out_8;
            arith_out_col_out_8_d2 <=  arith_out_col_out_8_d1;
            arith_out_col_out_8_d3 <=  arith_out_col_out_8_d2;
            arith_out_col_out_8_d4 <=  arith_out_col_out_8_d3;
            arith_out_col_out_8_d5 <=  arith_out_col_out_8_d4;
            arith_out_col_out_8_d6 <=  arith_out_col_out_8_d5;
            arith_out_col_out_8_d7 <=  arith_out_col_out_8_d6;
            arith_out_col_out_8_d8 <=  arith_out_col_out_8_d7;
            arith_out_col_out_8_d9 <=  arith_out_col_out_8_d8;
            arith_out_col_out_8_d10 <=  arith_out_col_out_8_d9;
            arith_out_col_out_8_d11 <=  arith_out_col_out_8_d10;
            arith_out_col_out_8_d12 <=  arith_out_col_out_8_d11;
            arith_out_col_out_8_d13 <=  arith_out_col_out_8_d12;
            arith_out_col_out_8_d14 <=  arith_out_col_out_8_d13;
            arith_out_col_out_8_d15 <=  arith_out_col_out_8_d14;
            arith_out_col_out_8_d16 <=  arith_out_col_out_8_d15;
            arith_out_col_out_8_d17 <=  arith_out_col_out_8_d16;
            arith_out_col_out_8_d18 <=  arith_out_col_out_8_d17;
            arith_out_col_out_8_d19 <=  arith_out_col_out_8_d18;
            arith_out_col_out_8_d20 <=  arith_out_col_out_8_d19;
            arith_out_col_out_8_d21 <=  arith_out_col_out_8_d20;
            arith_out_col_out_8_d22 <=  arith_out_col_out_8_d21;
            arith_out_col_out_9_d1 <=  arith_out_col_out_9;
            arith_out_col_out_9_d2 <=  arith_out_col_out_9_d1;
            arith_out_col_out_9_d3 <=  arith_out_col_out_9_d2;
            arith_out_col_out_9_d4 <=  arith_out_col_out_9_d3;
            arith_out_col_out_9_d5 <=  arith_out_col_out_9_d4;
            arith_out_col_out_9_d6 <=  arith_out_col_out_9_d5;
            arith_out_col_out_9_d7 <=  arith_out_col_out_9_d6;
            arith_out_col_out_9_d8 <=  arith_out_col_out_9_d7;
            arith_out_col_out_9_d9 <=  arith_out_col_out_9_d8;
            arith_out_col_out_9_d10 <=  arith_out_col_out_9_d9;
            arith_out_col_out_9_d11 <=  arith_out_col_out_9_d10;
            arith_out_col_out_9_d12 <=  arith_out_col_out_9_d11;
            arith_out_col_out_9_d13 <=  arith_out_col_out_9_d12;
            arith_out_col_out_9_d14 <=  arith_out_col_out_9_d13;
            arith_out_col_out_9_d15 <=  arith_out_col_out_9_d14;
            arith_out_col_out_9_d16 <=  arith_out_col_out_9_d15;
            arith_out_col_out_9_d17 <=  arith_out_col_out_9_d16;
            arith_out_col_out_9_d18 <=  arith_out_col_out_9_d17;
            arith_out_col_out_9_d19 <=  arith_out_col_out_9_d18;
            arith_out_col_out_9_d20 <=  arith_out_col_out_9_d19;
            arith_out_col_out_9_d21 <=  arith_out_col_out_9_d20;
            arith_out_col_out_10_d1 <=  arith_out_col_out_10;
            arith_out_col_out_10_d2 <=  arith_out_col_out_10_d1;
            arith_out_col_out_10_d3 <=  arith_out_col_out_10_d2;
            arith_out_col_out_10_d4 <=  arith_out_col_out_10_d3;
            arith_out_col_out_10_d5 <=  arith_out_col_out_10_d4;
            arith_out_col_out_10_d6 <=  arith_out_col_out_10_d5;
            arith_out_col_out_10_d7 <=  arith_out_col_out_10_d6;
            arith_out_col_out_10_d8 <=  arith_out_col_out_10_d7;
            arith_out_col_out_10_d9 <=  arith_out_col_out_10_d8;
            arith_out_col_out_10_d10 <=  arith_out_col_out_10_d9;
            arith_out_col_out_10_d11 <=  arith_out_col_out_10_d10;
            arith_out_col_out_10_d12 <=  arith_out_col_out_10_d11;
            arith_out_col_out_10_d13 <=  arith_out_col_out_10_d12;
            arith_out_col_out_10_d14 <=  arith_out_col_out_10_d13;
            arith_out_col_out_10_d15 <=  arith_out_col_out_10_d14;
            arith_out_col_out_10_d16 <=  arith_out_col_out_10_d15;
            arith_out_col_out_10_d17 <=  arith_out_col_out_10_d16;
            arith_out_col_out_10_d18 <=  arith_out_col_out_10_d17;
            arith_out_col_out_10_d19 <=  arith_out_col_out_10_d18;
            arith_out_col_out_10_d20 <=  arith_out_col_out_10_d19;
            arith_out_col_out_11_d1 <=  arith_out_col_out_11;
            arith_out_col_out_11_d2 <=  arith_out_col_out_11_d1;
            arith_out_col_out_11_d3 <=  arith_out_col_out_11_d2;
            arith_out_col_out_11_d4 <=  arith_out_col_out_11_d3;
            arith_out_col_out_11_d5 <=  arith_out_col_out_11_d4;
            arith_out_col_out_11_d6 <=  arith_out_col_out_11_d5;
            arith_out_col_out_11_d7 <=  arith_out_col_out_11_d6;
            arith_out_col_out_11_d8 <=  arith_out_col_out_11_d7;
            arith_out_col_out_11_d9 <=  arith_out_col_out_11_d8;
            arith_out_col_out_11_d10 <=  arith_out_col_out_11_d9;
            arith_out_col_out_11_d11 <=  arith_out_col_out_11_d10;
            arith_out_col_out_11_d12 <=  arith_out_col_out_11_d11;
            arith_out_col_out_11_d13 <=  arith_out_col_out_11_d12;
            arith_out_col_out_11_d14 <=  arith_out_col_out_11_d13;
            arith_out_col_out_11_d15 <=  arith_out_col_out_11_d14;
            arith_out_col_out_11_d16 <=  arith_out_col_out_11_d15;
            arith_out_col_out_11_d17 <=  arith_out_col_out_11_d16;
            arith_out_col_out_11_d18 <=  arith_out_col_out_11_d17;
            arith_out_col_out_11_d19 <=  arith_out_col_out_11_d18;
            arith_out_col_out_12_d1 <=  arith_out_col_out_12;
            arith_out_col_out_12_d2 <=  arith_out_col_out_12_d1;
            arith_out_col_out_12_d3 <=  arith_out_col_out_12_d2;
            arith_out_col_out_12_d4 <=  arith_out_col_out_12_d3;
            arith_out_col_out_12_d5 <=  arith_out_col_out_12_d4;
            arith_out_col_out_12_d6 <=  arith_out_col_out_12_d5;
            arith_out_col_out_12_d7 <=  arith_out_col_out_12_d6;
            arith_out_col_out_12_d8 <=  arith_out_col_out_12_d7;
            arith_out_col_out_12_d9 <=  arith_out_col_out_12_d8;
            arith_out_col_out_12_d10 <=  arith_out_col_out_12_d9;
            arith_out_col_out_12_d11 <=  arith_out_col_out_12_d10;
            arith_out_col_out_12_d12 <=  arith_out_col_out_12_d11;
            arith_out_col_out_12_d13 <=  arith_out_col_out_12_d12;
            arith_out_col_out_12_d14 <=  arith_out_col_out_12_d13;
            arith_out_col_out_12_d15 <=  arith_out_col_out_12_d14;
            arith_out_col_out_12_d16 <=  arith_out_col_out_12_d15;
            arith_out_col_out_12_d17 <=  arith_out_col_out_12_d16;
            arith_out_col_out_12_d18 <=  arith_out_col_out_12_d17;
            arith_out_col_out_13_d1 <=  arith_out_col_out_13;
            arith_out_col_out_13_d2 <=  arith_out_col_out_13_d1;
            arith_out_col_out_13_d3 <=  arith_out_col_out_13_d2;
            arith_out_col_out_13_d4 <=  arith_out_col_out_13_d3;
            arith_out_col_out_13_d5 <=  arith_out_col_out_13_d4;
            arith_out_col_out_13_d6 <=  arith_out_col_out_13_d5;
            arith_out_col_out_13_d7 <=  arith_out_col_out_13_d6;
            arith_out_col_out_13_d8 <=  arith_out_col_out_13_d7;
            arith_out_col_out_13_d9 <=  arith_out_col_out_13_d8;
            arith_out_col_out_13_d10 <=  arith_out_col_out_13_d9;
            arith_out_col_out_13_d11 <=  arith_out_col_out_13_d10;
            arith_out_col_out_13_d12 <=  arith_out_col_out_13_d11;
            arith_out_col_out_13_d13 <=  arith_out_col_out_13_d12;
            arith_out_col_out_13_d14 <=  arith_out_col_out_13_d13;
            arith_out_col_out_13_d15 <=  arith_out_col_out_13_d14;
            arith_out_col_out_13_d16 <=  arith_out_col_out_13_d15;
            arith_out_col_out_13_d17 <=  arith_out_col_out_13_d16;
            arith_out_col_out_14_d1 <=  arith_out_col_out_14;
            arith_out_col_out_14_d2 <=  arith_out_col_out_14_d1;
            arith_out_col_out_14_d3 <=  arith_out_col_out_14_d2;
            arith_out_col_out_14_d4 <=  arith_out_col_out_14_d3;
            arith_out_col_out_14_d5 <=  arith_out_col_out_14_d4;
            arith_out_col_out_14_d6 <=  arith_out_col_out_14_d5;
            arith_out_col_out_14_d7 <=  arith_out_col_out_14_d6;
            arith_out_col_out_14_d8 <=  arith_out_col_out_14_d7;
            arith_out_col_out_14_d9 <=  arith_out_col_out_14_d8;
            arith_out_col_out_14_d10 <=  arith_out_col_out_14_d9;
            arith_out_col_out_14_d11 <=  arith_out_col_out_14_d10;
            arith_out_col_out_14_d12 <=  arith_out_col_out_14_d11;
            arith_out_col_out_14_d13 <=  arith_out_col_out_14_d12;
            arith_out_col_out_14_d14 <=  arith_out_col_out_14_d13;
            arith_out_col_out_14_d15 <=  arith_out_col_out_14_d14;
            arith_out_col_out_14_d16 <=  arith_out_col_out_14_d15;
            arith_out_col_out_15_d1 <=  arith_out_col_out_15;
            arith_out_col_out_15_d2 <=  arith_out_col_out_15_d1;
            arith_out_col_out_15_d3 <=  arith_out_col_out_15_d2;
            arith_out_col_out_15_d4 <=  arith_out_col_out_15_d3;
            arith_out_col_out_15_d5 <=  arith_out_col_out_15_d4;
            arith_out_col_out_15_d6 <=  arith_out_col_out_15_d5;
            arith_out_col_out_15_d7 <=  arith_out_col_out_15_d6;
            arith_out_col_out_15_d8 <=  arith_out_col_out_15_d7;
            arith_out_col_out_15_d9 <=  arith_out_col_out_15_d8;
            arith_out_col_out_15_d10 <=  arith_out_col_out_15_d9;
            arith_out_col_out_15_d11 <=  arith_out_col_out_15_d10;
            arith_out_col_out_15_d12 <=  arith_out_col_out_15_d11;
            arith_out_col_out_15_d13 <=  arith_out_col_out_15_d12;
            arith_out_col_out_15_d14 <=  arith_out_col_out_15_d13;
            arith_out_col_out_15_d15 <=  arith_out_col_out_15_d14;
            arith_out_col_out_16_d1 <=  arith_out_col_out_16;
            arith_out_col_out_16_d2 <=  arith_out_col_out_16_d1;
            arith_out_col_out_16_d3 <=  arith_out_col_out_16_d2;
            arith_out_col_out_16_d4 <=  arith_out_col_out_16_d3;
            arith_out_col_out_16_d5 <=  arith_out_col_out_16_d4;
            arith_out_col_out_16_d6 <=  arith_out_col_out_16_d5;
            arith_out_col_out_16_d7 <=  arith_out_col_out_16_d6;
            arith_out_col_out_16_d8 <=  arith_out_col_out_16_d7;
            arith_out_col_out_16_d9 <=  arith_out_col_out_16_d8;
            arith_out_col_out_16_d10 <=  arith_out_col_out_16_d9;
            arith_out_col_out_16_d11 <=  arith_out_col_out_16_d10;
            arith_out_col_out_16_d12 <=  arith_out_col_out_16_d11;
            arith_out_col_out_16_d13 <=  arith_out_col_out_16_d12;
            arith_out_col_out_16_d14 <=  arith_out_col_out_16_d13;
            arith_out_col_out_17_d1 <=  arith_out_col_out_17;
            arith_out_col_out_17_d2 <=  arith_out_col_out_17_d1;
            arith_out_col_out_17_d3 <=  arith_out_col_out_17_d2;
            arith_out_col_out_17_d4 <=  arith_out_col_out_17_d3;
            arith_out_col_out_17_d5 <=  arith_out_col_out_17_d4;
            arith_out_col_out_17_d6 <=  arith_out_col_out_17_d5;
            arith_out_col_out_17_d7 <=  arith_out_col_out_17_d6;
            arith_out_col_out_17_d8 <=  arith_out_col_out_17_d7;
            arith_out_col_out_17_d9 <=  arith_out_col_out_17_d8;
            arith_out_col_out_17_d10 <=  arith_out_col_out_17_d9;
            arith_out_col_out_17_d11 <=  arith_out_col_out_17_d10;
            arith_out_col_out_17_d12 <=  arith_out_col_out_17_d11;
            arith_out_col_out_17_d13 <=  arith_out_col_out_17_d12;
            arith_out_col_out_18_d1 <=  arith_out_col_out_18;
            arith_out_col_out_18_d2 <=  arith_out_col_out_18_d1;
            arith_out_col_out_18_d3 <=  arith_out_col_out_18_d2;
            arith_out_col_out_18_d4 <=  arith_out_col_out_18_d3;
            arith_out_col_out_18_d5 <=  arith_out_col_out_18_d4;
            arith_out_col_out_18_d6 <=  arith_out_col_out_18_d5;
            arith_out_col_out_18_d7 <=  arith_out_col_out_18_d6;
            arith_out_col_out_18_d8 <=  arith_out_col_out_18_d7;
            arith_out_col_out_18_d9 <=  arith_out_col_out_18_d8;
            arith_out_col_out_18_d10 <=  arith_out_col_out_18_d9;
            arith_out_col_out_18_d11 <=  arith_out_col_out_18_d10;
            arith_out_col_out_18_d12 <=  arith_out_col_out_18_d11;
            arith_out_col_out_19_d1 <=  arith_out_col_out_19;
            arith_out_col_out_19_d2 <=  arith_out_col_out_19_d1;
            arith_out_col_out_19_d3 <=  arith_out_col_out_19_d2;
            arith_out_col_out_19_d4 <=  arith_out_col_out_19_d3;
            arith_out_col_out_19_d5 <=  arith_out_col_out_19_d4;
            arith_out_col_out_19_d6 <=  arith_out_col_out_19_d5;
            arith_out_col_out_19_d7 <=  arith_out_col_out_19_d6;
            arith_out_col_out_19_d8 <=  arith_out_col_out_19_d7;
            arith_out_col_out_19_d9 <=  arith_out_col_out_19_d8;
            arith_out_col_out_19_d10 <=  arith_out_col_out_19_d9;
            arith_out_col_out_19_d11 <=  arith_out_col_out_19_d10;
            arith_out_col_out_20_d1 <=  arith_out_col_out_20;
            arith_out_col_out_20_d2 <=  arith_out_col_out_20_d1;
            arith_out_col_out_20_d3 <=  arith_out_col_out_20_d2;
            arith_out_col_out_20_d4 <=  arith_out_col_out_20_d3;
            arith_out_col_out_20_d5 <=  arith_out_col_out_20_d4;
            arith_out_col_out_20_d6 <=  arith_out_col_out_20_d5;
            arith_out_col_out_20_d7 <=  arith_out_col_out_20_d6;
            arith_out_col_out_20_d8 <=  arith_out_col_out_20_d7;
            arith_out_col_out_20_d9 <=  arith_out_col_out_20_d8;
            arith_out_col_out_20_d10 <=  arith_out_col_out_20_d9;
            arith_out_col_out_21_d1 <=  arith_out_col_out_21;
            arith_out_col_out_21_d2 <=  arith_out_col_out_21_d1;
            arith_out_col_out_21_d3 <=  arith_out_col_out_21_d2;
            arith_out_col_out_21_d4 <=  arith_out_col_out_21_d3;
            arith_out_col_out_21_d5 <=  arith_out_col_out_21_d4;
            arith_out_col_out_21_d6 <=  arith_out_col_out_21_d5;
            arith_out_col_out_21_d7 <=  arith_out_col_out_21_d6;
            arith_out_col_out_21_d8 <=  arith_out_col_out_21_d7;
            arith_out_col_out_21_d9 <=  arith_out_col_out_21_d8;
            arith_out_col_out_22_d1 <=  arith_out_col_out_22;
            arith_out_col_out_22_d2 <=  arith_out_col_out_22_d1;
            arith_out_col_out_22_d3 <=  arith_out_col_out_22_d2;
            arith_out_col_out_22_d4 <=  arith_out_col_out_22_d3;
            arith_out_col_out_22_d5 <=  arith_out_col_out_22_d4;
            arith_out_col_out_22_d6 <=  arith_out_col_out_22_d5;
            arith_out_col_out_22_d7 <=  arith_out_col_out_22_d6;
            arith_out_col_out_22_d8 <=  arith_out_col_out_22_d7;
            arith_out_col_out_23_d1 <=  arith_out_col_out_23;
            arith_out_col_out_23_d2 <=  arith_out_col_out_23_d1;
            arith_out_col_out_23_d3 <=  arith_out_col_out_23_d2;
            arith_out_col_out_23_d4 <=  arith_out_col_out_23_d3;
            arith_out_col_out_23_d5 <=  arith_out_col_out_23_d4;
            arith_out_col_out_23_d6 <=  arith_out_col_out_23_d5;
            arith_out_col_out_23_d7 <=  arith_out_col_out_23_d6;
            arith_out_col_out_24_d1 <=  arith_out_col_out_24;
            arith_out_col_out_24_d2 <=  arith_out_col_out_24_d1;
            arith_out_col_out_24_d3 <=  arith_out_col_out_24_d2;
            arith_out_col_out_24_d4 <=  arith_out_col_out_24_d3;
            arith_out_col_out_24_d5 <=  arith_out_col_out_24_d4;
            arith_out_col_out_24_d6 <=  arith_out_col_out_24_d5;
            arith_out_col_out_25_d1 <=  arith_out_col_out_25;
            arith_out_col_out_25_d2 <=  arith_out_col_out_25_d1;
            arith_out_col_out_25_d3 <=  arith_out_col_out_25_d2;
            arith_out_col_out_25_d4 <=  arith_out_col_out_25_d3;
            arith_out_col_out_25_d5 <=  arith_out_col_out_25_d4;
            arith_out_col_out_26_d1 <=  arith_out_col_out_26;
            arith_out_col_out_26_d2 <=  arith_out_col_out_26_d1;
            arith_out_col_out_26_d3 <=  arith_out_col_out_26_d2;
            arith_out_col_out_26_d4 <=  arith_out_col_out_26_d3;
            arith_out_col_out_27_d1 <=  arith_out_col_out_27;
            arith_out_col_out_27_d2 <=  arith_out_col_out_27_d1;
            arith_out_col_out_27_d3 <=  arith_out_col_out_27_d2;
            arith_out_col_out_28_d1 <=  arith_out_col_out_28;
            arith_out_col_out_28_d2 <=  arith_out_col_out_28_d1;
            arith_out_col_out_29_d1 <=  arith_out_col_out_29;
         end if;
      end process;
------------ Delay depending on row index incoming dense arithmetic ------------
   arith_in_row_0 <= rowsA(3 downto 0);
   arith_in_row_0_q0 <= arith_in_row_0;
   arith_in_row_1 <= rowsA(7 downto 4);
   arith_in_row_1_q1 <= arith_in_row_1_d1;
   arith_in_row_2 <= rowsA(11 downto 8);
   arith_in_row_2_q2 <= arith_in_row_2_d2;
   arith_in_row_3 <= rowsA(15 downto 12);
   arith_in_row_3_q3 <= arith_in_row_3_d3;
   arith_in_row_4 <= rowsA(19 downto 16);
   arith_in_row_4_q4 <= arith_in_row_4_d4;
   arith_in_row_5 <= rowsA(23 downto 20);
   arith_in_row_5_q5 <= arith_in_row_5_d5;
   arith_in_row_6 <= rowsA(27 downto 24);
   arith_in_row_6_q6 <= arith_in_row_6_d6;
   arith_in_row_7 <= rowsA(31 downto 28);
   arith_in_row_7_q7 <= arith_in_row_7_d7;
   arith_in_row_8 <= rowsA(35 downto 32);
   arith_in_row_8_q8 <= arith_in_row_8_d8;
   arith_in_row_9 <= rowsA(39 downto 36);
   arith_in_row_9_q9 <= arith_in_row_9_d9;
   arith_in_row_10 <= rowsA(43 downto 40);
   arith_in_row_10_q10 <= arith_in_row_10_d10;
   arith_in_row_11 <= rowsA(47 downto 44);
   arith_in_row_11_q11 <= arith_in_row_11_d11;
   arith_in_row_12 <= rowsA(51 downto 48);
   arith_in_row_12_q12 <= arith_in_row_12_d12;
   arith_in_row_13 <= rowsA(55 downto 52);
   arith_in_row_13_q13 <= arith_in_row_13_d13;
   arith_in_row_14 <= rowsA(59 downto 56);
   arith_in_row_14_q14 <= arith_in_row_14_d14;
   arith_in_row_15 <= rowsA(63 downto 60);
   arith_in_row_15_q15 <= arith_in_row_15_d15;
   arith_in_row_16 <= rowsA(67 downto 64);
   arith_in_row_16_q16 <= arith_in_row_16_d16;
   arith_in_row_17 <= rowsA(71 downto 68);
   arith_in_row_17_q17 <= arith_in_row_17_d17;
   arith_in_row_18 <= rowsA(75 downto 72);
   arith_in_row_18_q18 <= arith_in_row_18_d18;
   arith_in_row_19 <= rowsA(79 downto 76);
   arith_in_row_19_q19 <= arith_in_row_19_d19;
   arith_in_row_20 <= rowsA(83 downto 80);
   arith_in_row_20_q20 <= arith_in_row_20_d20;
   arith_in_row_21 <= rowsA(87 downto 84);
   arith_in_row_21_q21 <= arith_in_row_21_d21;
   arith_in_row_22 <= rowsA(91 downto 88);
   arith_in_row_22_q22 <= arith_in_row_22_d22;
   arith_in_row_23 <= rowsA(95 downto 92);
   arith_in_row_23_q23 <= arith_in_row_23_d23;
   arith_in_row_24 <= rowsA(99 downto 96);
   arith_in_row_24_q24 <= arith_in_row_24_d24;
   arith_in_row_25 <= rowsA(103 downto 100);
   arith_in_row_25_q25 <= arith_in_row_25_d25;
   arith_in_row_26 <= rowsA(107 downto 104);
   arith_in_row_26_q26 <= arith_in_row_26_d26;
   arith_in_row_27 <= rowsA(111 downto 108);
   arith_in_row_27_q27 <= arith_in_row_27_d27;
   arith_in_row_28 <= rowsA(115 downto 112);
   arith_in_row_28_q28 <= arith_in_row_28_d28;
   arith_in_row_29 <= rowsA(119 downto 116);
   arith_in_row_29_q29 <= arith_in_row_29_d29;
   arith_in_row_30 <= rowsA(123 downto 120);
   arith_in_row_30_q30 <= arith_in_row_30_d30;
   arith_in_row_31 <= rowsA(127 downto 124);
   arith_in_row_31_q31 <= arith_in_row_31_d31;

------------ Delay depending on col index incoming dense arithmetic ------------
   arith_in_col_0 <= colsB(3 downto 0);
   arith_in_col_0_q0 <= arith_in_col_0;
   arith_in_col_1 <= colsB(7 downto 4);
   arith_in_col_1_q1 <= arith_in_col_1_d1;
   arith_in_col_2 <= colsB(11 downto 8);
   arith_in_col_2_q2 <= arith_in_col_2_d2;
   arith_in_col_3 <= colsB(15 downto 12);
   arith_in_col_3_q3 <= arith_in_col_3_d3;
   arith_in_col_4 <= colsB(19 downto 16);
   arith_in_col_4_q4 <= arith_in_col_4_d4;
   arith_in_col_5 <= colsB(23 downto 20);
   arith_in_col_5_q5 <= arith_in_col_5_d5;
   arith_in_col_6 <= colsB(27 downto 24);
   arith_in_col_6_q6 <= arith_in_col_6_d6;
   arith_in_col_7 <= colsB(31 downto 28);
   arith_in_col_7_q7 <= arith_in_col_7_d7;
   arith_in_col_8 <= colsB(35 downto 32);
   arith_in_col_8_q8 <= arith_in_col_8_d8;
   arith_in_col_9 <= colsB(39 downto 36);
   arith_in_col_9_q9 <= arith_in_col_9_d9;
   arith_in_col_10 <= colsB(43 downto 40);
   arith_in_col_10_q10 <= arith_in_col_10_d10;
   arith_in_col_11 <= colsB(47 downto 44);
   arith_in_col_11_q11 <= arith_in_col_11_d11;
   arith_in_col_12 <= colsB(51 downto 48);
   arith_in_col_12_q12 <= arith_in_col_12_d12;
   arith_in_col_13 <= colsB(55 downto 52);
   arith_in_col_13_q13 <= arith_in_col_13_d13;
   arith_in_col_14 <= colsB(59 downto 56);
   arith_in_col_14_q14 <= arith_in_col_14_d14;
   arith_in_col_15 <= colsB(63 downto 60);
   arith_in_col_15_q15 <= arith_in_col_15_d15;
   arith_in_col_16 <= colsB(67 downto 64);
   arith_in_col_16_q16 <= arith_in_col_16_d16;
   arith_in_col_17 <= colsB(71 downto 68);
   arith_in_col_17_q17 <= arith_in_col_17_d17;
   arith_in_col_18 <= colsB(75 downto 72);
   arith_in_col_18_q18 <= arith_in_col_18_d18;
   arith_in_col_19 <= colsB(79 downto 76);
   arith_in_col_19_q19 <= arith_in_col_19_d19;
   arith_in_col_20 <= colsB(83 downto 80);
   arith_in_col_20_q20 <= arith_in_col_20_d20;
   arith_in_col_21 <= colsB(87 downto 84);
   arith_in_col_21_q21 <= arith_in_col_21_d21;
   arith_in_col_22 <= colsB(91 downto 88);
   arith_in_col_22_q22 <= arith_in_col_22_d22;
   arith_in_col_23 <= colsB(95 downto 92);
   arith_in_col_23_q23 <= arith_in_col_23_d23;
   arith_in_col_24 <= colsB(99 downto 96);
   arith_in_col_24_q24 <= arith_in_col_24_d24;
   arith_in_col_25 <= colsB(103 downto 100);
   arith_in_col_25_q25 <= arith_in_col_25_d25;
   arith_in_col_26 <= colsB(107 downto 104);
   arith_in_col_26_q26 <= arith_in_col_26_d26;
   arith_in_col_27 <= colsB(111 downto 108);
   arith_in_col_27_q27 <= arith_in_col_27_d27;
   arith_in_col_28 <= colsB(115 downto 112);
   arith_in_col_28_q28 <= arith_in_col_28_d28;
   arith_in_col_29 <= colsB(119 downto 116);
   arith_in_col_29_q29 <= arith_in_col_29_d29;
   arith_in_col_30 <= colsB(123 downto 120);
   arith_in_col_30_q30 <= arith_in_col_30_d30;

--------------- Delay SOB/EOB with Arith_to_S3 delay to feed SAK ---------------
   SOB_select <= SOB;
   SOB_q0 <= SOB_select;
   EOB_select <= EOB;
   EOB_q0 <= EOB_select;

--------------- Delay outgoing arithmetic depending on col index ---------------
   arith_out_col_out_0 <= LAICPT2_to_arith(3 downto 0);
   arith_out_col_out_0_q30 <= arith_out_col_out_0_d30;
   arith_out_col_out_1 <= LAICPT2_to_arith(7 downto 4);
   arith_out_col_out_1_q29 <= arith_out_col_out_1_d29;
   arith_out_col_out_2 <= LAICPT2_to_arith(11 downto 8);
   arith_out_col_out_2_q28 <= arith_out_col_out_2_d28;
   arith_out_col_out_3 <= LAICPT2_to_arith(15 downto 12);
   arith_out_col_out_3_q27 <= arith_out_col_out_3_d27;
   arith_out_col_out_4 <= LAICPT2_to_arith(19 downto 16);
   arith_out_col_out_4_q26 <= arith_out_col_out_4_d26;
   arith_out_col_out_5 <= LAICPT2_to_arith(23 downto 20);
   arith_out_col_out_5_q25 <= arith_out_col_out_5_d25;
   arith_out_col_out_6 <= LAICPT2_to_arith(27 downto 24);
   arith_out_col_out_6_q24 <= arith_out_col_out_6_d24;
   arith_out_col_out_7 <= LAICPT2_to_arith(31 downto 28);
   arith_out_col_out_7_q23 <= arith_out_col_out_7_d23;
   arith_out_col_out_8 <= LAICPT2_to_arith(35 downto 32);
   arith_out_col_out_8_q22 <= arith_out_col_out_8_d22;
   arith_out_col_out_9 <= LAICPT2_to_arith(39 downto 36);
   arith_out_col_out_9_q21 <= arith_out_col_out_9_d21;
   arith_out_col_out_10 <= LAICPT2_to_arith(43 downto 40);
   arith_out_col_out_10_q20 <= arith_out_col_out_10_d20;
   arith_out_col_out_11 <= LAICPT2_to_arith(47 downto 44);
   arith_out_col_out_11_q19 <= arith_out_col_out_11_d19;
   arith_out_col_out_12 <= LAICPT2_to_arith(51 downto 48);
   arith_out_col_out_12_q18 <= arith_out_col_out_12_d18;
   arith_out_col_out_13 <= LAICPT2_to_arith(55 downto 52);
   arith_out_col_out_13_q17 <= arith_out_col_out_13_d17;
   arith_out_col_out_14 <= LAICPT2_to_arith(59 downto 56);
   arith_out_col_out_14_q16 <= arith_out_col_out_14_d16;
   arith_out_col_out_15 <= LAICPT2_to_arith(63 downto 60);
   arith_out_col_out_15_q15 <= arith_out_col_out_15_d15;
   arith_out_col_out_16 <= LAICPT2_to_arith(67 downto 64);
   arith_out_col_out_16_q14 <= arith_out_col_out_16_d14;
   arith_out_col_out_17 <= LAICPT2_to_arith(71 downto 68);
   arith_out_col_out_17_q13 <= arith_out_col_out_17_d13;
   arith_out_col_out_18 <= LAICPT2_to_arith(75 downto 72);
   arith_out_col_out_18_q12 <= arith_out_col_out_18_d12;
   arith_out_col_out_19 <= LAICPT2_to_arith(79 downto 76);
   arith_out_col_out_19_q11 <= arith_out_col_out_19_d11;
   arith_out_col_out_20 <= LAICPT2_to_arith(83 downto 80);
   arith_out_col_out_20_q10 <= arith_out_col_out_20_d10;
   arith_out_col_out_21 <= LAICPT2_to_arith(87 downto 84);
   arith_out_col_out_21_q9 <= arith_out_col_out_21_d9;
   arith_out_col_out_22 <= LAICPT2_to_arith(91 downto 88);
   arith_out_col_out_22_q8 <= arith_out_col_out_22_d8;
   arith_out_col_out_23 <= LAICPT2_to_arith(95 downto 92);
   arith_out_col_out_23_q7 <= arith_out_col_out_23_d7;
   arith_out_col_out_24 <= LAICPT2_to_arith(99 downto 96);
   arith_out_col_out_24_q6 <= arith_out_col_out_24_d6;
   arith_out_col_out_25 <= LAICPT2_to_arith(103 downto 100);
   arith_out_col_out_25_q5 <= arith_out_col_out_25_d5;
   arith_out_col_out_26 <= LAICPT2_to_arith(107 downto 104);
   arith_out_col_out_26_q4 <= arith_out_col_out_26_d4;
   arith_out_col_out_27 <= LAICPT2_to_arith(111 downto 108);
   arith_out_col_out_27_q3 <= arith_out_col_out_27_d3;
   arith_out_col_out_28 <= LAICPT2_to_arith(115 downto 112);
   arith_out_col_out_28_q2 <= arith_out_col_out_28_d2;
   arith_out_col_out_29 <= LAICPT2_to_arith(119 downto 116);
   arith_out_col_out_29_q1 <= arith_out_col_out_29_d1;
   arith_out_col_out_30 <= LAICPT2_to_arith(123 downto 120);
   arith_out_col_out_30_q0 <= arith_out_col_out_30;

---------------- Generate Arith_to_S3 for rows and connect them ----------------
   rows_i_arith(0) <= arith_in_row_0_q0;
   rows_i_arith(1) <= arith_in_row_1_q1;
   rows_i_arith(2) <= arith_in_row_2_q2;
   rows_i_arith(3) <= arith_in_row_3_q3;
   rows_i_arith(4) <= arith_in_row_4_q4;
   rows_i_arith(5) <= arith_in_row_5_q5;
   rows_i_arith(6) <= arith_in_row_6_q6;
   rows_i_arith(7) <= arith_in_row_7_q7;
   rows_i_arith(8) <= arith_in_row_8_q8;
   rows_i_arith(9) <= arith_in_row_9_q9;
   rows_i_arith(10) <= arith_in_row_10_q10;
   rows_i_arith(11) <= arith_in_row_11_q11;
   rows_i_arith(12) <= arith_in_row_12_q12;
   rows_i_arith(13) <= arith_in_row_13_q13;
   rows_i_arith(14) <= arith_in_row_14_q14;
   rows_i_arith(15) <= arith_in_row_15_q15;
   rows_i_arith(16) <= arith_in_row_16_q16;
   rows_i_arith(17) <= arith_in_row_17_q17;
   rows_i_arith(18) <= arith_in_row_18_q18;
   rows_i_arith(19) <= arith_in_row_19_q19;
   rows_i_arith(20) <= arith_in_row_20_q20;
   rows_i_arith(21) <= arith_in_row_21_q21;
   rows_i_arith(22) <= arith_in_row_22_q22;
   rows_i_arith(23) <= arith_in_row_23_q23;
   rows_i_arith(24) <= arith_in_row_24_q24;
   rows_i_arith(25) <= arith_in_row_25_q25;
   rows_i_arith(26) <= arith_in_row_26_q26;
   rows_i_arith(27) <= arith_in_row_27_q27;
   rows_i_arith(28) <= arith_in_row_28_q28;
   rows_i_arith(29) <= arith_in_row_29_q29;
   rows_i_arith(30) <= arith_in_row_30_q30;
   rows_i_arith(31) <= arith_in_row_31_q31;
   rows_a2s3: for II in 0 to 31 generate
      a2s3_i: Arith_to_S3
         port map ( clk => clk,
                    arith_i => rows_i_arith(II),
                    s3_o => rows_i_s3(((II+1)*7)-1 downto II*7));
   end generate;

---------------- Generate Arith_to_S3 for cols and connect them ----------------
   cols_j_arith(0) <= arith_in_col_0_q0;
   cols_j_arith(1) <= arith_in_col_1_q1;
   cols_j_arith(2) <= arith_in_col_2_q2;
   cols_j_arith(3) <= arith_in_col_3_q3;
   cols_j_arith(4) <= arith_in_col_4_q4;
   cols_j_arith(5) <= arith_in_col_5_q5;
   cols_j_arith(6) <= arith_in_col_6_q6;
   cols_j_arith(7) <= arith_in_col_7_q7;
   cols_j_arith(8) <= arith_in_col_8_q8;
   cols_j_arith(9) <= arith_in_col_9_q9;
   cols_j_arith(10) <= arith_in_col_10_q10;
   cols_j_arith(11) <= arith_in_col_11_q11;
   cols_j_arith(12) <= arith_in_col_12_q12;
   cols_j_arith(13) <= arith_in_col_13_q13;
   cols_j_arith(14) <= arith_in_col_14_q14;
   cols_j_arith(15) <= arith_in_col_15_q15;
   cols_j_arith(16) <= arith_in_col_16_q16;
   cols_j_arith(17) <= arith_in_col_17_q17;
   cols_j_arith(18) <= arith_in_col_18_q18;
   cols_j_arith(19) <= arith_in_col_19_q19;
   cols_j_arith(20) <= arith_in_col_20_q20;
   cols_j_arith(21) <= arith_in_col_21_q21;
   cols_j_arith(22) <= arith_in_col_22_q22;
   cols_j_arith(23) <= arith_in_col_23_q23;
   cols_j_arith(24) <= arith_in_col_24_q24;
   cols_j_arith(25) <= arith_in_col_25_q25;
   cols_j_arith(26) <= arith_in_col_26_q26;
   cols_j_arith(27) <= arith_in_col_27_q27;
   cols_j_arith(28) <= arith_in_col_28_q28;
   cols_j_arith(29) <= arith_in_col_29_q29;
   cols_j_arith(30) <= arith_in_col_30_q30;
   cols_a2s3: for JJ in 0 to 30 generate
      a2s3_j: Arith_to_S3
         port map ( clk => clk,
                    arith_i => cols_j_arith(JJ),
                    s3_o => cols_j_s3(((JJ+1)*7)-1 downto JJ*7));
   end generate;

-------------------- Instantiate the Systolic Array Kernel --------------------
   sak: SystolicArrayKernel
      port map ( clk => clk,
                 rst => rst,
                 rowsA => rows_i_s3,
                 colsB => cols_j_s3,
                 SOB => SOB_q0,
                 EOB => EOB_q0,
                 EOB_Q_o => EOB_Q_o,
                 colsC => colsC_LAICPT2 );

-------------------------- Generate LAICPT2_to_arith --------------------------
   cols_l2a: for JJ in 0 to 30 generate
      l2a_i: l2a
         port map ( clk => clk,
                    A => colsC_LAICPT2(((JJ+1)*15)-1-1-0 downto JJ*15),
                    isNaN => colsC_LAICPT2(((JJ+1)*15)- 1),
                    arith_o => LAICPT2_to_arith(((JJ+1)*4)-1 downto JJ*4));
   end generate;

-------- Connect outgoing delayed dense arith words to colsC output bus --------
   colsC(3 downto 0) <= arith_out_col_out_0_q30;
   colsC(7 downto 4) <= arith_out_col_out_1_q29;
   colsC(11 downto 8) <= arith_out_col_out_2_q28;
   colsC(15 downto 12) <= arith_out_col_out_3_q27;
   colsC(19 downto 16) <= arith_out_col_out_4_q26;
   colsC(23 downto 20) <= arith_out_col_out_5_q25;
   colsC(27 downto 24) <= arith_out_col_out_6_q24;
   colsC(31 downto 28) <= arith_out_col_out_7_q23;
   colsC(35 downto 32) <= arith_out_col_out_8_q22;
   colsC(39 downto 36) <= arith_out_col_out_9_q21;
   colsC(43 downto 40) <= arith_out_col_out_10_q20;
   colsC(47 downto 44) <= arith_out_col_out_11_q19;
   colsC(51 downto 48) <= arith_out_col_out_12_q18;
   colsC(55 downto 52) <= arith_out_col_out_13_q17;
   colsC(59 downto 56) <= arith_out_col_out_14_q16;
   colsC(63 downto 60) <= arith_out_col_out_15_q15;
   colsC(67 downto 64) <= arith_out_col_out_16_q14;
   colsC(71 downto 68) <= arith_out_col_out_17_q13;
   colsC(75 downto 72) <= arith_out_col_out_18_q12;
   colsC(79 downto 76) <= arith_out_col_out_19_q11;
   colsC(83 downto 80) <= arith_out_col_out_20_q10;
   colsC(87 downto 84) <= arith_out_col_out_21_q9;
   colsC(91 downto 88) <= arith_out_col_out_22_q8;
   colsC(95 downto 92) <= arith_out_col_out_23_q7;
   colsC(99 downto 96) <= arith_out_col_out_24_q6;
   colsC(103 downto 100) <= arith_out_col_out_25_q5;
   colsC(107 downto 104) <= arith_out_col_out_26_q4;
   colsC(111 downto 108) <= arith_out_col_out_27_q3;
   colsC(115 downto 112) <= arith_out_col_out_28_q2;
   colsC(119 downto 116) <= arith_out_col_out_29_q1;
   colsC(123 downto 120) <= arith_out_col_out_30_q0;

end architecture;

