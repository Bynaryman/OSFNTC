--------------------------------------------------------------------------------
--                            MultTable_F200_uid40
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid40 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid40 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_F200_uid45
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid45 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid45 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_F200_uid50
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid50 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid50 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_F200_uid55
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid55 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid55 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_F200_uid60
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid60 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid60 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_F200_uid65
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid65 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid65 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_F200_uid70
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid70 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid70 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_F200_uid75
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid75 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid75 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_F200_uid80
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid80 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid80 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_F200_uid85
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid85 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid85 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_F200_uid90
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid90 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid90 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                            MultTable_F200_uid95
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid95 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid95 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid110
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid110 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid110 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid115
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid115 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid115 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid120
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid120 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid120 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid125
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid125 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid125 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid130
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid130 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid130 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid135
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid135 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid135 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid140
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid140 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid140 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid145
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid145 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid145 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid150
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid150 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid150 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid155
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid155 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid155 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid160
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid160 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid160 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid165
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid165 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid165 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid180
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid180 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid180 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid185
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid185 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid185 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid190
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid190 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid190 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid195
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid195 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid195 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid200
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid200 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid200 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid205
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid205 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid205 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid210
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid210 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid210 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid215
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid215 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid215 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid220
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid220 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid220 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid225
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid225 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid225 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid230
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid230 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid230 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid235
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid235 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid235 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid240
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid240 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid240 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid245
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid245 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid245 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                        Compressor_23_3_F200_uid249
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_F200_uid249 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_F200_uid249 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                         Compressor_3_2_F200_uid257
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_F200_uid257 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_F200_uid257 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                        Compressor_14_3_F200_uid271
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_F200_uid271 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_F200_uid271 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                         Compressor_6_3_F200_uid305
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_F200_uid305 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_F200_uid305 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid823
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid823 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid823 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid828
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid828 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid828 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid833
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid833 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid833 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid838
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid838 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid838 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid843
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid843 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid843 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid848
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid848 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid848 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid853
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid853 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid853 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid858
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid858 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid858 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid863
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid863 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid863 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid868
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid868 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid868 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid873
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid873 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid873 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid878
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid878 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid878 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid893
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid893 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid893 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid898
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid898 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid898 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid903
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid903 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid903 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid908
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid908 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid908 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid913
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid913 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid913 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid918
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid918 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid918 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid923
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid923 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid923 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid928
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid928 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid928 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid933
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid933 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid933 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid938
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid938 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid938 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid943
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid943 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid943 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid948
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid948 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid948 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid963
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid963 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid963 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid968
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid968 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid968 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid973
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid973 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid973 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid978
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid978 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid978 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid983
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid983 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid983 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid988
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid988 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid988 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid993
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid993 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid993 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid998
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid998 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid998 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid1003
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid1003 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid1003 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid1008
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid1008 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid1008 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid1013
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid1013 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid1013 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid1018
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid1018 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid1018 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid1023
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid1023 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid1023 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                           MultTable_F200_uid1028
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_F200_uid1028 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_F200_uid1028 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                        Compressor_23_3_F200_uid1032
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_F200_uid1032 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_F200_uid1032 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                        Compressor_3_2_F200_uid1040
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_F200_uid1040 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_F200_uid1040 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                        Compressor_14_3_F200_uid1054
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_F200_uid1054 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_F200_uid1054 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                        Compressor_6_3_F200_uid1088
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_F200_uid1088 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_F200_uid1088 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                                Arith_to_S3
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: BSC / UPC - Ledoux Louis
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: arith_i
-- Output signals: S3_o

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Arith_to_S3 is
    port (clk : in std_logic;
          arith_i : in  std_logic_vector(63 downto 0);
          S3_o : out  std_logic_vector(65 downto 0)   );
end entity;

architecture arch of Arith_to_S3 is
signal sign :  std_logic;
signal exponent :  std_logic_vector(10 downto 0);
signal fraction :  std_logic_vector(51 downto 0);
signal isNaN :  std_logic;
signal isExpSubnormalZero :  std_logic;
signal implicit :  std_logic;
signal final_scale :  std_logic_vector(10 downto 0);
begin
   sign <= arith_i(63);
   exponent <= arith_i(62 downto 52);
   fraction <= arith_i(51 downto 0);
   isNaN <= '1' when exponent="11111111111" else '0';
   isExpSubnormalZero <= '1' when exponent="00000000000" else '0';
   implicit <= not(isExpSubnormalZero);
   final_scale<= "00000000001" when isExpSubnormalZero= '1' else  exponent;
   S3_o <= isNaN & sign & implicit & fraction & final_scale;
end architecture;

--------------------------------------------------------------------------------
--            LZOCShifterSticky_100_to_54_counting_128_F200_uid784
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: I OZb
-- Output signals: Count O Sticky

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZOCShifterSticky_100_to_54_counting_128_F200_uid784 is
    port (clk : in std_logic;
          I : in  std_logic_vector(99 downto 0);
          OZb : in  std_logic;
          Count : out  std_logic_vector(6 downto 0);
          O : out  std_logic_vector(53 downto 0);
          Sticky : out  std_logic   );
end entity;

architecture arch of LZOCShifterSticky_100_to_54_counting_128_F200_uid784 is
signal level7 :  std_logic_vector(99 downto 0);
signal sozb, sozb_d1, sozb_d2 :  std_logic;
signal sticky7 :  std_logic;
signal count6, count6_d1, count6_d2 :  std_logic;
signal level6 :  std_logic_vector(99 downto 0);
signal sticky_high_6 :  std_logic;
signal sticky_low_6 :  std_logic;
signal sticky6 :  std_logic;
signal count5, count5_d1, count5_d2 :  std_logic;
signal level5, level5_d1 :  std_logic_vector(84 downto 0);
signal sticky_high_5 :  std_logic;
signal sticky_low_5 :  std_logic;
signal sticky5, sticky5_d1 :  std_logic;
signal count4, count4_d1 :  std_logic;
signal level4 :  std_logic_vector(68 downto 0);
signal sticky_high_4, sticky_high_4_d1 :  std_logic;
signal sticky_low_4, sticky_low_4_d1 :  std_logic;
signal sticky4 :  std_logic;
signal count3, count3_d1 :  std_logic;
signal level3 :  std_logic_vector(60 downto 0);
signal sticky_high_3 :  std_logic;
signal sticky_low_3, sticky_low_3_d1 :  std_logic;
signal sticky3 :  std_logic;
signal count2, count2_d1 :  std_logic;
signal level2, level2_d1 :  std_logic_vector(56 downto 0);
signal sticky_high_2 :  std_logic;
signal sticky_low_2, sticky_low_2_d1 :  std_logic;
signal sticky2, sticky2_d1 :  std_logic;
signal count1, count1_d1 :  std_logic;
signal level1 :  std_logic_vector(54 downto 0);
signal sticky_high_1, sticky_high_1_d1 :  std_logic;
signal sticky_low_1, sticky_low_1_d1, sticky_low_1_d2 :  std_logic;
signal sticky1 :  std_logic;
signal count0 :  std_logic;
signal level0 :  std_logic_vector(53 downto 0);
signal sticky_high_0 :  std_logic;
signal sticky_low_0, sticky_low_0_d1, sticky_low_0_d2 :  std_logic;
signal sticky0 :  std_logic;
signal sCount :  std_logic_vector(6 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sozb_d1 <=  sozb;
            sozb_d2 <=  sozb_d1;
            count6_d1 <=  count6;
            count6_d2 <=  count6_d1;
            count5_d1 <=  count5;
            count5_d2 <=  count5_d1;
            level5_d1 <=  level5;
            sticky5_d1 <=  sticky5;
            count4_d1 <=  count4;
            sticky_high_4_d1 <=  sticky_high_4;
            sticky_low_4_d1 <=  sticky_low_4;
            count3_d1 <=  count3;
            sticky_low_3_d1 <=  sticky_low_3;
            count2_d1 <=  count2;
            level2_d1 <=  level2;
            sticky_low_2_d1 <=  sticky_low_2;
            sticky2_d1 <=  sticky2;
            count1_d1 <=  count1;
            sticky_high_1_d1 <=  sticky_high_1;
            sticky_low_1_d1 <=  sticky_low_1;
            sticky_low_1_d2 <=  sticky_low_1_d1;
            sticky_low_0_d1 <=  sticky_low_0;
            sticky_low_0_d2 <=  sticky_low_0_d1;
         end if;
      end process;
   level7 <= I ;
   sozb<= OZb;
   sticky7 <= '0' ;
   count6<= '1' when level7(99 downto 36) = (99 downto 36=>sozb) else '0';
   level6<= level7(99 downto 0) when count6='0' else level7(35 downto 0) & (63 downto 0 => '0');
   sticky_high_6<= '0';
   sticky_low_6<= '0';
   sticky6<= sticky7 or sticky_high_6 when count6='0' else sticky7 or sticky_low_6;

   count5<= '1' when level6(99 downto 68) = (99 downto 68=>sozb) else '0';
   level5<= level6(99 downto 15) when count5='0' else level6(67 downto 0) & (16 downto 0 => '0');
   sticky_high_5<= '0'when level6(14 downto 0) = CONV_STD_LOGIC_VECTOR(0,15) else '1';
   sticky_low_5<= '0';
   sticky5<= sticky6 or sticky_high_5 when count5='0' else sticky6 or sticky_low_5;

   count4<= '1' when level5_d1(84 downto 69) = (84 downto 69=>sozb_d1) else '0';
   level4<= level5_d1(84 downto 16) when count4='0' else level5_d1(68 downto 0);
   sticky_high_4<= '0'when level5(15 downto 0) = CONV_STD_LOGIC_VECTOR(0,16) else '1';
   sticky_low_4<= '0';
   sticky4<= sticky5_d1 or sticky_high_4_d1 when count4='0' else sticky5_d1 or sticky_low_4_d1;

   count3<= '1' when level4(68 downto 61) = (68 downto 61=>sozb_d1) else '0';
   level3<= level4(68 downto 8) when count3='0' else level4(60 downto 0);
   sticky_high_3<= '0'when level4(7 downto 0) = CONV_STD_LOGIC_VECTOR(0,8) else '1';
   sticky_low_3<= '0';
   sticky3<= sticky4 or sticky_high_3 when count3='0' else sticky4 or sticky_low_3_d1;

   count2<= '1' when level3(60 downto 57) = (60 downto 57=>sozb_d1) else '0';
   level2<= level3(60 downto 4) when count2='0' else level3(56 downto 0);
   sticky_high_2<= '0'when level3(3 downto 0) = CONV_STD_LOGIC_VECTOR(0,4) else '1';
   sticky_low_2<= '0';
   sticky2<= sticky3 or sticky_high_2 when count2='0' else sticky3 or sticky_low_2_d1;

   count1<= '1' when level2(56 downto 55) = (56 downto 55=>sozb_d1) else '0';
   level1<= level2_d1(56 downto 2) when count1_d1='0' else level2_d1(54 downto 0);
   sticky_high_1<= '0'when level2(1 downto 0) = CONV_STD_LOGIC_VECTOR(0,2) else '1';
   sticky_low_1<= '0';
   sticky1<= sticky2_d1 or sticky_high_1_d1 when count1_d1='0' else sticky2_d1 or sticky_low_1_d2;

   count0<= '1' when level1(54 downto 54) = (54 downto 54=>sozb_d2) else '0';
   level0<= level1(54 downto 1) when count0='0' else level1(53 downto 0);
   sticky_high_0<= '0'when level1(0 downto 0) = CONV_STD_LOGIC_VECTOR(0,1) else '1';
   sticky_low_0<= '0';
   sticky0<= sticky1 or sticky_high_0 when count0='0' else sticky1 or sticky_low_0_d2;

   O <= level0;
   sCount <= count6_d2 & count5_d2 & count4_d1 & count3_d1 & count2_d1 & count1_d1 & count0;
   Count <= sCount;
   Sticky <= sticky0;
end architecture;

--------------------------------------------------------------------------------
--                                    l2a
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Ledoux Louis - BSC / UPC
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: A isNaN
-- Output signals: arith_o

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity l2a is
    port (clk : in std_logic;
          A : in  std_logic_vector(99 downto 0);
          isNaN : in  std_logic;
          arith_o : out  std_logic_vector(63 downto 0)   );
end entity;

architecture arch of l2a is
   component LZOCShifterSticky_100_to_54_counting_128_F200_uid784 is
      port ( clk : in std_logic;
             I : in  std_logic_vector(99 downto 0);
             OZb : in  std_logic;
             Count : out  std_logic_vector(6 downto 0);
             O : out  std_logic_vector(53 downto 0);
             Sticky : out  std_logic   );
   end component;

signal rippled_carry, rippled_carry_d1, rippled_carry_d2 :  std_logic_vector(99 downto 0);
signal count_bit :  std_logic;
signal count_lzoc_o :  std_logic_vector(6 downto 0);
signal frac_lzoc_o :  std_logic_vector(53 downto 0);
signal sticky_lzoc_o :  std_logic;
signal unbiased_exp :  std_logic_vector(6 downto 0);
signal bias, bias_d1, bias_d2 :  std_logic_vector(10 downto 0);
signal biased_exp :  std_logic_vector(10 downto 0);
signal not_frac_lzoc :  std_logic_vector(53 downto 0);
signal unrounded_frac :  std_logic_vector(53 downto 0);
signal G :  std_logic;
signal R :  std_logic;
signal S :  std_logic;
signal round_up :  std_logic;
signal rounded_frac :  std_logic_vector(53 downto 0);
signal post_round_ovf :  std_logic;
signal post_rounding_exp :  std_logic_vector(11 downto 0);
signal nan_out :  std_logic;
signal is_zero :  std_logic;
signal final_exp :  std_logic_vector(10 downto 0);
signal isNaN_d1, isNaN_d2 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            rippled_carry_d1 <=  rippled_carry;
            rippled_carry_d2 <=  rippled_carry_d1;
            bias_d1 <=  bias;
            bias_d2 <=  bias_d1;
            isNaN_d1 <=  isNaN;
            isNaN_d2 <=  isNaN_d1;
         end if;
      end process;

   rippled_carry <= A;

--------------- Count 0/1 while shifting and sticky computation ---------------
   count_bit <= rippled_carry(99);
   lzoc_inst: LZOCShifterSticky_100_to_54_counting_128_F200_uid784
      port map ( clk  => clk,
                 I => rippled_carry,
                 OZb => count_bit,
                 Count => count_lzoc_o,
                 O => frac_lzoc_o,
                 Sticky => sticky_lzoc_o);

----------- Compute unbiased exponent from msb weigth and lzoc count -----------
   unbiased_exp <= CONV_STD_LOGIC_VECTOR(49,7) - (count_lzoc_o);
   bias <= CONV_STD_LOGIC_VECTOR(1023,11);
   biased_exp <= bias_d2 + ((10 downto 7 => unbiased_exp(6)) & unbiased_exp);

-------------------------- Convert in sign magnitude --------------------------
   not_frac_lzoc <=  frac_lzoc_o xor (53 downto 0 => rippled_carry_d2(99));
   unrounded_frac <= "0" & not_frac_lzoc(52 downto 0) + rippled_carry_d2(99);

---- G and R should be taken from lzoc adding one size more frac lzoc width ----
------------------------------- GRS rounding up -------------------------------
   G <= unrounded_frac(1);
   R <= unrounded_frac(0);
   S <= sticky_lzoc_o;
   round_up <= G and (R or S);
   rounded_frac <= unrounded_frac + round_up;
   post_round_ovf <= rounded_frac(53);

------------------------- post rounding scale handling -------------------------
   post_rounding_exp <= ("0" & biased_exp) + (rounded_frac(53));
   nan_out <= post_rounding_exp(11) or isNaN_d2;
is_zero <= count_lzoc_o(6) when rounded_frac="000000000000000000000000000000000000000000000000000000" else '0';
   final_exp <= post_rounding_exp(10 downto 0) when nan_out = '0' else "11111111111";
   arith_o <= (rippled_carry_d2(99) & final_exp(10 downto 0) & rounded_frac(52 downto 1)) when is_zero = '0' else "0000000000000000000000000000000000000000000000000000000000000000";
end architecture;

--------------------------------------------------------------------------------
--                         DSPBlock_17x24_F200_uid795
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_F200_uid795 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_F200_uid795 is
signal Mint :  std_logic_vector(40 downto 0);
signal M :  std_logic_vector(40 downto 0);
signal Rtmp :  std_logic_vector(40 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(40 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                         DSPBlock_17x24_F200_uid797
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_F200_uid797 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_F200_uid797 is
signal Mint :  std_logic_vector(40 downto 0);
signal M :  std_logic_vector(40 downto 0);
signal Rtmp :  std_logic_vector(40 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(40 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                         DSPBlock_17x24_F200_uid799
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_F200_uid799 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_F200_uid799 is
signal Mint :  std_logic_vector(40 downto 0);
signal M :  std_logic_vector(40 downto 0);
signal Rtmp :  std_logic_vector(40 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(40 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                         DSPBlock_2x24_F200_uid801
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_2x24_F200_uid801 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(25 downto 0)   );
end entity;

architecture arch of DSPBlock_2x24_F200_uid801 is
signal Mint :  std_logic_vector(25 downto 0);
signal M :  std_logic_vector(25 downto 0);
signal Rtmp :  std_logic_vector(25 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(25 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                         DSPBlock_17x24_F200_uid803
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_F200_uid803 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_F200_uid803 is
signal Mint :  std_logic_vector(40 downto 0);
signal M :  std_logic_vector(40 downto 0);
signal Rtmp :  std_logic_vector(40 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(40 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                         DSPBlock_17x24_F200_uid805
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_F200_uid805 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_F200_uid805 is
signal Mint :  std_logic_vector(40 downto 0);
signal M :  std_logic_vector(40 downto 0);
signal Rtmp :  std_logic_vector(40 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(40 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                         DSPBlock_17x24_F200_uid807
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_F200_uid807 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_F200_uid807 is
signal Mint :  std_logic_vector(40 downto 0);
signal M :  std_logic_vector(40 downto 0);
signal Rtmp :  std_logic_vector(40 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(40 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                         DSPBlock_2x24_F200_uid809
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_2x24_F200_uid809 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(25 downto 0)   );
end entity;

architecture arch of DSPBlock_2x24_F200_uid809 is
signal Mint :  std_logic_vector(25 downto 0);
signal M :  std_logic_vector(25 downto 0);
signal Rtmp :  std_logic_vector(25 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(25 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_1x1_F200_uid811
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_F200_uid811 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_F200_uid811 is
signal replicated :  std_logic_vector(0 downto 0);
signal prod :  std_logic_vector(0 downto 0);
begin
   replicated <= (0 downto 0 => X(0));
   prod <= Y and replicated;
   R <= prod;
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_4x1_F200_uid813
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_F200_uid813 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_F200_uid813 is
signal replicated :  std_logic_vector(3 downto 0);
signal prod :  std_logic_vector(3 downto 0);
begin
   replicated <= (3 downto 0 => Y(0));
   prod <= X and replicated;
   R <= prod;
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_4x1_F200_uid815
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_F200_uid815 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_F200_uid815 is
signal replicated :  std_logic_vector(3 downto 0);
signal prod :  std_logic_vector(3 downto 0);
begin
   replicated <= (3 downto 0 => Y(0));
   prod <= X and replicated;
   R <= prod;
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_4x1_F200_uid817
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_F200_uid817 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_F200_uid817 is
signal replicated :  std_logic_vector(3 downto 0);
signal prod :  std_logic_vector(3 downto 0);
begin
   replicated <= (3 downto 0 => Y(0));
   prod <= X and replicated;
   R <= prod;
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_4x1_F200_uid819
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_F200_uid819 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_F200_uid819 is
signal replicated :  std_logic_vector(3 downto 0);
signal prod :  std_logic_vector(3 downto 0);
begin
   replicated <= (3 downto 0 => Y(0));
   prod <= X and replicated;
   R <= prod;
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_2x2_F200_uid821
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_F200_uid821 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_F200_uid821 is
   component MultTable_F200_uid823 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(3 downto 0);
signal Y1 :  std_logic_vector(3 downto 0);
signal Y1_copy824 :  std_logic_vector(3 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid823
      port map ( X => Xtable,
                 Y => Y1_copy824);
   Y1 <= Y1_copy824; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid826
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid826 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid826 is
   component MultTable_F200_uid828 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy829 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid828
      port map ( X => Xtable,
                 Y => Y1_copy829);
   Y1 <= Y1_copy829; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid831
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid831 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid831 is
   component MultTable_F200_uid833 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy834 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid833
      port map ( X => Xtable,
                 Y => Y1_copy834);
   Y1 <= Y1_copy834; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid836
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid836 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid836 is
   component MultTable_F200_uid838 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy839 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid838
      port map ( X => Xtable,
                 Y => Y1_copy839);
   Y1 <= Y1_copy839; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid841
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid841 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid841 is
   component MultTable_F200_uid843 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy844 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid843
      port map ( X => Xtable,
                 Y => Y1_copy844);
   Y1 <= Y1_copy844; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid846
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid846 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid846 is
   component MultTable_F200_uid848 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy849 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid848
      port map ( X => Xtable,
                 Y => Y1_copy849);
   Y1 <= Y1_copy849; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_2x2_F200_uid851
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_F200_uid851 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_F200_uid851 is
   component MultTable_F200_uid853 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(3 downto 0);
signal Y1 :  std_logic_vector(3 downto 0);
signal Y1_copy854 :  std_logic_vector(3 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid853
      port map ( X => Xtable,
                 Y => Y1_copy854);
   Y1 <= Y1_copy854; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid856
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid856 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid856 is
   component MultTable_F200_uid858 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy859 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid858
      port map ( X => Xtable,
                 Y => Y1_copy859);
   Y1 <= Y1_copy859; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid861
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid861 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid861 is
   component MultTable_F200_uid863 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy864 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid863
      port map ( X => Xtable,
                 Y => Y1_copy864);
   Y1 <= Y1_copy864; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid866
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid866 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid866 is
   component MultTable_F200_uid868 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy869 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid868
      port map ( X => Xtable,
                 Y => Y1_copy869);
   Y1 <= Y1_copy869; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid871
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid871 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid871 is
   component MultTable_F200_uid873 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy874 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid873
      port map ( X => Xtable,
                 Y => Y1_copy874);
   Y1 <= Y1_copy874; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid876
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid876 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid876 is
   component MultTable_F200_uid878 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy879 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid878
      port map ( X => Xtable,
                 Y => Y1_copy879);
   Y1 <= Y1_copy879; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_1x1_F200_uid881
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_F200_uid881 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_F200_uid881 is
signal replicated :  std_logic_vector(0 downto 0);
signal prod :  std_logic_vector(0 downto 0);
begin
   replicated <= (0 downto 0 => X(0));
   prod <= Y and replicated;
   R <= prod;
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_4x1_F200_uid883
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_F200_uid883 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_F200_uid883 is
signal replicated :  std_logic_vector(3 downto 0);
signal prod :  std_logic_vector(3 downto 0);
begin
   replicated <= (3 downto 0 => Y(0));
   prod <= X and replicated;
   R <= prod;
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_4x1_F200_uid885
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_F200_uid885 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_F200_uid885 is
signal replicated :  std_logic_vector(3 downto 0);
signal prod :  std_logic_vector(3 downto 0);
begin
   replicated <= (3 downto 0 => Y(0));
   prod <= X and replicated;
   R <= prod;
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_4x1_F200_uid887
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_F200_uid887 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_F200_uid887 is
signal replicated :  std_logic_vector(3 downto 0);
signal prod :  std_logic_vector(3 downto 0);
begin
   replicated <= (3 downto 0 => Y(0));
   prod <= X and replicated;
   R <= prod;
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_4x1_F200_uid889
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_F200_uid889 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_F200_uid889 is
signal replicated :  std_logic_vector(3 downto 0);
signal prod :  std_logic_vector(3 downto 0);
begin
   replicated <= (3 downto 0 => Y(0));
   prod <= X and replicated;
   R <= prod;
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_2x2_F200_uid891
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_F200_uid891 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_F200_uid891 is
   component MultTable_F200_uid893 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(3 downto 0);
signal Y1 :  std_logic_vector(3 downto 0);
signal Y1_copy894 :  std_logic_vector(3 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid893
      port map ( X => Xtable,
                 Y => Y1_copy894);
   Y1 <= Y1_copy894; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid896
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid896 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid896 is
   component MultTable_F200_uid898 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy899 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid898
      port map ( X => Xtable,
                 Y => Y1_copy899);
   Y1 <= Y1_copy899; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid901
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid901 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid901 is
   component MultTable_F200_uid903 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy904 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid903
      port map ( X => Xtable,
                 Y => Y1_copy904);
   Y1 <= Y1_copy904; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid906
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid906 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid906 is
   component MultTable_F200_uid908 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy909 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid908
      port map ( X => Xtable,
                 Y => Y1_copy909);
   Y1 <= Y1_copy909; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid911
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid911 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid911 is
   component MultTable_F200_uid913 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy914 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid913
      port map ( X => Xtable,
                 Y => Y1_copy914);
   Y1 <= Y1_copy914; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid916
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid916 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid916 is
   component MultTable_F200_uid918 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy919 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid918
      port map ( X => Xtable,
                 Y => Y1_copy919);
   Y1 <= Y1_copy919; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_2x2_F200_uid921
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_F200_uid921 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_F200_uid921 is
   component MultTable_F200_uid923 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(3 downto 0);
signal Y1 :  std_logic_vector(3 downto 0);
signal Y1_copy924 :  std_logic_vector(3 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid923
      port map ( X => Xtable,
                 Y => Y1_copy924);
   Y1 <= Y1_copy924; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid926
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid926 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid926 is
   component MultTable_F200_uid928 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy929 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid928
      port map ( X => Xtable,
                 Y => Y1_copy929);
   Y1 <= Y1_copy929; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid931
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid931 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid931 is
   component MultTable_F200_uid933 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy934 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid933
      port map ( X => Xtable,
                 Y => Y1_copy934);
   Y1 <= Y1_copy934; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid936
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid936 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid936 is
   component MultTable_F200_uid938 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy939 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid938
      port map ( X => Xtable,
                 Y => Y1_copy939);
   Y1 <= Y1_copy939; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid941
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid941 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid941 is
   component MultTable_F200_uid943 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy944 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid943
      port map ( X => Xtable,
                 Y => Y1_copy944);
   Y1 <= Y1_copy944; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid946
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid946 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid946 is
   component MultTable_F200_uid948 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy949 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid948
      port map ( X => Xtable,
                 Y => Y1_copy949);
   Y1 <= Y1_copy949; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_1x1_F200_uid951
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_F200_uid951 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_F200_uid951 is
signal replicated :  std_logic_vector(0 downto 0);
signal prod :  std_logic_vector(0 downto 0);
begin
   replicated <= (0 downto 0 => X(0));
   prod <= Y and replicated;
   R <= prod;
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_4x1_F200_uid953
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_F200_uid953 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_F200_uid953 is
signal replicated :  std_logic_vector(3 downto 0);
signal prod :  std_logic_vector(3 downto 0);
begin
   replicated <= (3 downto 0 => Y(0));
   prod <= X and replicated;
   R <= prod;
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_4x1_F200_uid955
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_F200_uid955 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_F200_uid955 is
signal replicated :  std_logic_vector(3 downto 0);
signal prod :  std_logic_vector(3 downto 0);
begin
   replicated <= (3 downto 0 => Y(0));
   prod <= X and replicated;
   R <= prod;
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_4x1_F200_uid957
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_F200_uid957 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_F200_uid957 is
signal replicated :  std_logic_vector(3 downto 0);
signal prod :  std_logic_vector(3 downto 0);
begin
   replicated <= (3 downto 0 => Y(0));
   prod <= X and replicated;
   R <= prod;
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_4x1_F200_uid959
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_F200_uid959 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_F200_uid959 is
signal replicated :  std_logic_vector(3 downto 0);
signal prod :  std_logic_vector(3 downto 0);
begin
   replicated <= (3 downto 0 => Y(0));
   prod <= X and replicated;
   R <= prod;
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_2x2_F200_uid961
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_F200_uid961 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_F200_uid961 is
   component MultTable_F200_uid963 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(3 downto 0);
signal Y1 :  std_logic_vector(3 downto 0);
signal Y1_copy964 :  std_logic_vector(3 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid963
      port map ( X => Xtable,
                 Y => Y1_copy964);
   Y1 <= Y1_copy964; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid966
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid966 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid966 is
   component MultTable_F200_uid968 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy969 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid968
      port map ( X => Xtable,
                 Y => Y1_copy969);
   Y1 <= Y1_copy969; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid971
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid971 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid971 is
   component MultTable_F200_uid973 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy974 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid973
      port map ( X => Xtable,
                 Y => Y1_copy974);
   Y1 <= Y1_copy974; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid976
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid976 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid976 is
   component MultTable_F200_uid978 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy979 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid978
      port map ( X => Xtable,
                 Y => Y1_copy979);
   Y1 <= Y1_copy979; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid981
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid981 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid981 is
   component MultTable_F200_uid983 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy984 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid983
      port map ( X => Xtable,
                 Y => Y1_copy984);
   Y1 <= Y1_copy984; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid986
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid986 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid986 is
   component MultTable_F200_uid988 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy989 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid988
      port map ( X => Xtable,
                 Y => Y1_copy989);
   Y1 <= Y1_copy989; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_2x2_F200_uid991
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_F200_uid991 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_F200_uid991 is
   component MultTable_F200_uid993 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(3 downto 0);
signal Y1 :  std_logic_vector(3 downto 0);
signal Y1_copy994 :  std_logic_vector(3 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid993
      port map ( X => Xtable,
                 Y => Y1_copy994);
   Y1 <= Y1_copy994; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiplierLUT_3x2_F200_uid996
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid996 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid996 is
   component MultTable_F200_uid998 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy999 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid998
      port map ( X => Xtable,
                 Y => Y1_copy999);
   Y1 <= Y1_copy999; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_F200_uid1001
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid1001 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid1001 is
   component MultTable_F200_uid1003 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy1004 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid1003
      port map ( X => Xtable,
                 Y => Y1_copy1004);
   Y1 <= Y1_copy1004; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_F200_uid1006
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid1006 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid1006 is
   component MultTable_F200_uid1008 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy1009 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid1008
      port map ( X => Xtable,
                 Y => Y1_copy1009);
   Y1 <= Y1_copy1009; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_F200_uid1011
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid1011 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid1011 is
   component MultTable_F200_uid1013 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy1014 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid1013
      port map ( X => Xtable,
                 Y => Y1_copy1014);
   Y1 <= Y1_copy1014; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_F200_uid1016
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_F200_uid1016 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_F200_uid1016 is
   component MultTable_F200_uid1018 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy1019 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid1018
      port map ( X => Xtable,
                 Y => Y1_copy1019);
   Y1 <= Y1_copy1019; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x2_F200_uid1021
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_F200_uid1021 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_F200_uid1021 is
   component MultTable_F200_uid1023 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(3 downto 0);
signal Y1 :  std_logic_vector(3 downto 0);
signal Y1_copy1024 :  std_logic_vector(3 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid1023
      port map ( X => Xtable,
                 Y => Y1_copy1024);
   Y1 <= Y1_copy1024; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_F200_uid1026
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_F200_uid1026 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_F200_uid1026 is
   component MultTable_F200_uid1028 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable :  std_logic_vector(4 downto 0);
signal Y1 :  std_logic_vector(4 downto 0);
signal Y1_copy1029 :  std_logic_vector(4 downto 0);
begin
Xtable <= Y & X;
   R <= Y1;
   TableMult: MultTable_F200_uid1028
      port map ( X => Xtable,
                 Y => Y1_copy1029);
   Y1 <= Y1_copy1029; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_82_F200_uid1560
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_82_F200_uid1560 is
    port (clk : in std_logic;
          X : in  std_logic_vector(81 downto 0);
          Y : in  std_logic_vector(81 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(81 downto 0)   );
end entity;

architecture arch of IntAdder_82_F200_uid1560 is
signal Rtmp :  std_logic_vector(81 downto 0);
begin
   Rtmp <= X + Y + Cin;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                         IntMultiplier_F200_uid791
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_F200_uid791 is
    port (clk : in std_logic;
          X : in  std_logic_vector(52 downto 0);
          Y : in  std_logic_vector(52 downto 0);
          R : out  std_logic_vector(105 downto 0)   );
end entity;

architecture arch of IntMultiplier_F200_uid791 is
   component DSPBlock_17x24_F200_uid795 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_F200_uid797 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_F200_uid799 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_2x24_F200_uid801 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(25 downto 0)   );
   end component;

   component DSPBlock_17x24_F200_uid803 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_F200_uid805 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_F200_uid807 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_2x24_F200_uid809 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(25 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_F200_uid811 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_F200_uid813 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_F200_uid815 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_F200_uid817 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_F200_uid819 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_F200_uid821 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid826 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid831 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid836 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid841 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid846 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_F200_uid851 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid856 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid861 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid866 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid871 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid876 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_F200_uid881 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_F200_uid883 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_F200_uid885 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_F200_uid887 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_F200_uid889 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_F200_uid891 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid896 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid901 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid906 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid911 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid916 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_F200_uid921 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid926 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid931 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid936 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid941 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid946 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_F200_uid951 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_F200_uid953 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_F200_uid955 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_F200_uid957 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_F200_uid959 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_F200_uid961 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid966 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid971 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid976 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid981 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid986 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_F200_uid991 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid996 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid1001 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid1006 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid1011 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_F200_uid1016 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_F200_uid1021 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_F200_uid1026 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_F200_uid1032 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_F200_uid1040 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component Compressor_14_3_F200_uid1054 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_6_3_F200_uid1088 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_82_F200_uid1560 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(81 downto 0);
             Y : in  std_logic_vector(81 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(81 downto 0)   );
   end component;

signal XX_m792 :  std_logic_vector(52 downto 0);
signal YY_m792 :  std_logic_vector(52 downto 0);
signal tile_0_X :  std_logic_vector(16 downto 0);
signal tile_0_Y :  std_logic_vector(23 downto 0);
signal tile_0_output :  std_logic_vector(40 downto 0);
signal tile_0_filtered_output :  std_logic_vector(40 downto 0);
signal bh793_w0_0 :  std_logic;
signal bh793_w1_0 :  std_logic;
signal bh793_w2_0 :  std_logic;
signal bh793_w3_0 :  std_logic;
signal bh793_w4_0 :  std_logic;
signal bh793_w5_0 :  std_logic;
signal bh793_w6_0 :  std_logic;
signal bh793_w7_0 :  std_logic;
signal bh793_w8_0 :  std_logic;
signal bh793_w9_0 :  std_logic;
signal bh793_w10_0 :  std_logic;
signal bh793_w11_0 :  std_logic;
signal bh793_w12_0 :  std_logic;
signal bh793_w13_0 :  std_logic;
signal bh793_w14_0 :  std_logic;
signal bh793_w15_0 :  std_logic;
signal bh793_w16_0 :  std_logic;
signal bh793_w17_0 :  std_logic;
signal bh793_w18_0 :  std_logic;
signal bh793_w19_0 :  std_logic;
signal bh793_w20_0 :  std_logic;
signal bh793_w21_0 :  std_logic;
signal bh793_w22_0 :  std_logic;
signal bh793_w23_0 :  std_logic;
signal bh793_w24_0 :  std_logic;
signal bh793_w25_0 :  std_logic;
signal bh793_w26_0 :  std_logic;
signal bh793_w27_0 :  std_logic;
signal bh793_w28_0 :  std_logic;
signal bh793_w29_0 :  std_logic;
signal bh793_w30_0 :  std_logic;
signal bh793_w31_0 :  std_logic;
signal bh793_w32_0 :  std_logic;
signal bh793_w33_0 :  std_logic;
signal bh793_w34_0 :  std_logic;
signal bh793_w35_0 :  std_logic;
signal bh793_w36_0 :  std_logic;
signal bh793_w37_0 :  std_logic;
signal bh793_w38_0 :  std_logic;
signal bh793_w39_0 :  std_logic;
signal bh793_w40_0 :  std_logic;
signal tile_1_X :  std_logic_vector(16 downto 0);
signal tile_1_Y :  std_logic_vector(23 downto 0);
signal tile_1_output :  std_logic_vector(40 downto 0);
signal tile_1_filtered_output :  std_logic_vector(40 downto 0);
signal bh793_w17_1 :  std_logic;
signal bh793_w18_1 :  std_logic;
signal bh793_w19_1 :  std_logic;
signal bh793_w20_1 :  std_logic;
signal bh793_w21_1 :  std_logic;
signal bh793_w22_1 :  std_logic;
signal bh793_w23_1 :  std_logic;
signal bh793_w24_1 :  std_logic;
signal bh793_w25_1 :  std_logic;
signal bh793_w26_1 :  std_logic;
signal bh793_w27_1 :  std_logic;
signal bh793_w28_1 :  std_logic;
signal bh793_w29_1 :  std_logic;
signal bh793_w30_1 :  std_logic;
signal bh793_w31_1 :  std_logic;
signal bh793_w32_1 :  std_logic;
signal bh793_w33_1 :  std_logic;
signal bh793_w34_1 :  std_logic;
signal bh793_w35_1 :  std_logic;
signal bh793_w36_1 :  std_logic;
signal bh793_w37_1 :  std_logic;
signal bh793_w38_1 :  std_logic;
signal bh793_w39_1 :  std_logic;
signal bh793_w40_1 :  std_logic;
signal bh793_w41_0 :  std_logic;
signal bh793_w42_0 :  std_logic;
signal bh793_w43_0 :  std_logic;
signal bh793_w44_0 :  std_logic;
signal bh793_w45_0 :  std_logic;
signal bh793_w46_0 :  std_logic;
signal bh793_w47_0 :  std_logic;
signal bh793_w48_0 :  std_logic;
signal bh793_w49_0 :  std_logic;
signal bh793_w50_0 :  std_logic;
signal bh793_w51_0 :  std_logic;
signal bh793_w52_0 :  std_logic;
signal bh793_w53_0 :  std_logic;
signal bh793_w54_0 :  std_logic;
signal bh793_w55_0 :  std_logic;
signal bh793_w56_0 :  std_logic;
signal bh793_w57_0 :  std_logic;
signal tile_2_X :  std_logic_vector(16 downto 0);
signal tile_2_Y :  std_logic_vector(23 downto 0);
signal tile_2_output :  std_logic_vector(40 downto 0);
signal tile_2_filtered_output :  std_logic_vector(40 downto 0);
signal bh793_w34_2 :  std_logic;
signal bh793_w35_2 :  std_logic;
signal bh793_w36_2 :  std_logic;
signal bh793_w37_2 :  std_logic;
signal bh793_w38_2 :  std_logic;
signal bh793_w39_2 :  std_logic;
signal bh793_w40_2 :  std_logic;
signal bh793_w41_1 :  std_logic;
signal bh793_w42_1 :  std_logic;
signal bh793_w43_1 :  std_logic;
signal bh793_w44_1 :  std_logic;
signal bh793_w45_1 :  std_logic;
signal bh793_w46_1 :  std_logic;
signal bh793_w47_1 :  std_logic;
signal bh793_w48_1 :  std_logic;
signal bh793_w49_1 :  std_logic;
signal bh793_w50_1 :  std_logic;
signal bh793_w51_1 :  std_logic;
signal bh793_w52_1 :  std_logic;
signal bh793_w53_1 :  std_logic;
signal bh793_w54_1 :  std_logic;
signal bh793_w55_1 :  std_logic;
signal bh793_w56_1 :  std_logic;
signal bh793_w57_1 :  std_logic;
signal bh793_w58_0 :  std_logic;
signal bh793_w59_0 :  std_logic;
signal bh793_w60_0 :  std_logic;
signal bh793_w61_0 :  std_logic;
signal bh793_w62_0 :  std_logic;
signal bh793_w63_0 :  std_logic;
signal bh793_w64_0 :  std_logic;
signal bh793_w65_0 :  std_logic;
signal bh793_w66_0 :  std_logic;
signal bh793_w67_0 :  std_logic;
signal bh793_w68_0 :  std_logic;
signal bh793_w69_0 :  std_logic;
signal bh793_w70_0 :  std_logic;
signal bh793_w71_0 :  std_logic;
signal bh793_w72_0 :  std_logic;
signal bh793_w73_0 :  std_logic;
signal bh793_w74_0 :  std_logic;
signal tile_3_X :  std_logic_vector(1 downto 0);
signal tile_3_Y :  std_logic_vector(23 downto 0);
signal tile_3_output :  std_logic_vector(25 downto 0);
signal tile_3_filtered_output :  std_logic_vector(25 downto 0);
signal bh793_w51_2 :  std_logic;
signal bh793_w52_2 :  std_logic;
signal bh793_w53_2 :  std_logic;
signal bh793_w54_2 :  std_logic;
signal bh793_w55_2 :  std_logic;
signal bh793_w56_2 :  std_logic;
signal bh793_w57_2 :  std_logic;
signal bh793_w58_1 :  std_logic;
signal bh793_w59_1 :  std_logic;
signal bh793_w60_1 :  std_logic;
signal bh793_w61_1 :  std_logic;
signal bh793_w62_1 :  std_logic;
signal bh793_w63_1 :  std_logic;
signal bh793_w64_1 :  std_logic;
signal bh793_w65_1 :  std_logic;
signal bh793_w66_1 :  std_logic;
signal bh793_w67_1 :  std_logic;
signal bh793_w68_1 :  std_logic;
signal bh793_w69_1 :  std_logic;
signal bh793_w70_1 :  std_logic;
signal bh793_w71_1 :  std_logic;
signal bh793_w72_1 :  std_logic;
signal bh793_w73_1 :  std_logic;
signal bh793_w74_1 :  std_logic;
signal bh793_w75_0 :  std_logic;
signal bh793_w76_0 :  std_logic;
signal tile_4_X :  std_logic_vector(16 downto 0);
signal tile_4_Y :  std_logic_vector(23 downto 0);
signal tile_4_output :  std_logic_vector(40 downto 0);
signal tile_4_filtered_output :  std_logic_vector(40 downto 0);
signal bh793_w24_2 :  std_logic;
signal bh793_w25_2 :  std_logic;
signal bh793_w26_2 :  std_logic;
signal bh793_w27_2 :  std_logic;
signal bh793_w28_2 :  std_logic;
signal bh793_w29_2 :  std_logic;
signal bh793_w30_2 :  std_logic;
signal bh793_w31_2 :  std_logic;
signal bh793_w32_2 :  std_logic;
signal bh793_w33_2 :  std_logic;
signal bh793_w34_3 :  std_logic;
signal bh793_w35_3 :  std_logic;
signal bh793_w36_3 :  std_logic;
signal bh793_w37_3 :  std_logic;
signal bh793_w38_3 :  std_logic;
signal bh793_w39_3 :  std_logic;
signal bh793_w40_3 :  std_logic;
signal bh793_w41_2 :  std_logic;
signal bh793_w42_2 :  std_logic;
signal bh793_w43_2 :  std_logic;
signal bh793_w44_2 :  std_logic;
signal bh793_w45_2 :  std_logic;
signal bh793_w46_2 :  std_logic;
signal bh793_w47_2 :  std_logic;
signal bh793_w48_2 :  std_logic;
signal bh793_w49_2 :  std_logic;
signal bh793_w50_2 :  std_logic;
signal bh793_w51_3 :  std_logic;
signal bh793_w52_3 :  std_logic;
signal bh793_w53_3 :  std_logic;
signal bh793_w54_3 :  std_logic;
signal bh793_w55_3 :  std_logic;
signal bh793_w56_3 :  std_logic;
signal bh793_w57_3 :  std_logic;
signal bh793_w58_2 :  std_logic;
signal bh793_w59_2 :  std_logic;
signal bh793_w60_2 :  std_logic;
signal bh793_w61_2 :  std_logic;
signal bh793_w62_2 :  std_logic;
signal bh793_w63_2 :  std_logic;
signal bh793_w64_2 :  std_logic;
signal tile_5_X :  std_logic_vector(16 downto 0);
signal tile_5_Y :  std_logic_vector(23 downto 0);
signal tile_5_output :  std_logic_vector(40 downto 0);
signal tile_5_filtered_output :  std_logic_vector(40 downto 0);
signal bh793_w41_3 :  std_logic;
signal bh793_w42_3 :  std_logic;
signal bh793_w43_3 :  std_logic;
signal bh793_w44_3 :  std_logic;
signal bh793_w45_3 :  std_logic;
signal bh793_w46_3 :  std_logic;
signal bh793_w47_3 :  std_logic;
signal bh793_w48_3 :  std_logic;
signal bh793_w49_3 :  std_logic;
signal bh793_w50_3 :  std_logic;
signal bh793_w51_4 :  std_logic;
signal bh793_w52_4 :  std_logic;
signal bh793_w53_4 :  std_logic;
signal bh793_w54_4 :  std_logic;
signal bh793_w55_4 :  std_logic;
signal bh793_w56_4 :  std_logic;
signal bh793_w57_4 :  std_logic;
signal bh793_w58_3 :  std_logic;
signal bh793_w59_3 :  std_logic;
signal bh793_w60_3 :  std_logic;
signal bh793_w61_3 :  std_logic;
signal bh793_w62_3 :  std_logic;
signal bh793_w63_3 :  std_logic;
signal bh793_w64_3 :  std_logic;
signal bh793_w65_2 :  std_logic;
signal bh793_w66_2 :  std_logic;
signal bh793_w67_2 :  std_logic;
signal bh793_w68_2 :  std_logic;
signal bh793_w69_2 :  std_logic;
signal bh793_w70_2 :  std_logic;
signal bh793_w71_2 :  std_logic;
signal bh793_w72_2 :  std_logic;
signal bh793_w73_2 :  std_logic;
signal bh793_w74_2 :  std_logic;
signal bh793_w75_1 :  std_logic;
signal bh793_w76_1 :  std_logic;
signal bh793_w77_0 :  std_logic;
signal bh793_w78_0 :  std_logic;
signal bh793_w79_0 :  std_logic;
signal bh793_w80_0 :  std_logic;
signal bh793_w81_0 :  std_logic;
signal tile_6_X :  std_logic_vector(16 downto 0);
signal tile_6_Y :  std_logic_vector(23 downto 0);
signal tile_6_output :  std_logic_vector(40 downto 0);
signal tile_6_filtered_output :  std_logic_vector(40 downto 0);
signal bh793_w58_4 :  std_logic;
signal bh793_w59_4 :  std_logic;
signal bh793_w60_4 :  std_logic;
signal bh793_w61_4 :  std_logic;
signal bh793_w62_4 :  std_logic;
signal bh793_w63_4 :  std_logic;
signal bh793_w64_4 :  std_logic;
signal bh793_w65_3 :  std_logic;
signal bh793_w66_3 :  std_logic;
signal bh793_w67_3 :  std_logic;
signal bh793_w68_3 :  std_logic;
signal bh793_w69_3 :  std_logic;
signal bh793_w70_3 :  std_logic;
signal bh793_w71_3 :  std_logic;
signal bh793_w72_3 :  std_logic;
signal bh793_w73_3 :  std_logic;
signal bh793_w74_3 :  std_logic;
signal bh793_w75_2 :  std_logic;
signal bh793_w76_2 :  std_logic;
signal bh793_w77_1 :  std_logic;
signal bh793_w78_1 :  std_logic;
signal bh793_w79_1 :  std_logic;
signal bh793_w80_1 :  std_logic;
signal bh793_w81_1 :  std_logic;
signal bh793_w82_0 :  std_logic;
signal bh793_w83_0 :  std_logic;
signal bh793_w84_0 :  std_logic;
signal bh793_w85_0 :  std_logic;
signal bh793_w86_0 :  std_logic;
signal bh793_w87_0 :  std_logic;
signal bh793_w88_0 :  std_logic;
signal bh793_w89_0 :  std_logic;
signal bh793_w90_0 :  std_logic;
signal bh793_w91_0 :  std_logic;
signal bh793_w92_0 :  std_logic;
signal bh793_w93_0 :  std_logic;
signal bh793_w94_0 :  std_logic;
signal bh793_w95_0 :  std_logic;
signal bh793_w96_0 :  std_logic;
signal bh793_w97_0 :  std_logic;
signal bh793_w98_0 :  std_logic;
signal tile_7_X :  std_logic_vector(1 downto 0);
signal tile_7_Y :  std_logic_vector(23 downto 0);
signal tile_7_output :  std_logic_vector(25 downto 0);
signal tile_7_filtered_output :  std_logic_vector(25 downto 0);
signal bh793_w75_3 :  std_logic;
signal bh793_w76_3 :  std_logic;
signal bh793_w77_2 :  std_logic;
signal bh793_w78_2 :  std_logic;
signal bh793_w79_2 :  std_logic;
signal bh793_w80_2 :  std_logic;
signal bh793_w81_2 :  std_logic;
signal bh793_w82_1 :  std_logic;
signal bh793_w83_1 :  std_logic;
signal bh793_w84_1 :  std_logic;
signal bh793_w85_1 :  std_logic;
signal bh793_w86_1 :  std_logic;
signal bh793_w87_1 :  std_logic;
signal bh793_w88_1 :  std_logic;
signal bh793_w89_1 :  std_logic;
signal bh793_w90_1 :  std_logic;
signal bh793_w91_1 :  std_logic;
signal bh793_w92_1 :  std_logic;
signal bh793_w93_1 :  std_logic;
signal bh793_w94_1 :  std_logic;
signal bh793_w95_1 :  std_logic;
signal bh793_w96_1 :  std_logic;
signal bh793_w97_1 :  std_logic;
signal bh793_w98_1 :  std_logic;
signal bh793_w99_0 :  std_logic;
signal bh793_w100_0 :  std_logic;
signal tile_8_X :  std_logic_vector(0 downto 0);
signal tile_8_Y :  std_logic_vector(0 downto 0);
signal tile_8_output :  std_logic_vector(0 downto 0);
signal tile_8_filtered_output :  std_logic_vector(0 downto 0);
signal bh793_w68_4 :  std_logic;
signal tile_9_X :  std_logic_vector(3 downto 0);
signal tile_9_Y :  std_logic_vector(0 downto 0);
signal tile_9_output :  std_logic_vector(3 downto 0);
signal tile_9_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w64_5 :  std_logic;
signal bh793_w65_4 :  std_logic;
signal bh793_w66_4 :  std_logic;
signal bh793_w67_4 :  std_logic;
signal tile_10_X :  std_logic_vector(3 downto 0);
signal tile_10_Y :  std_logic_vector(0 downto 0);
signal tile_10_output :  std_logic_vector(3 downto 0);
signal tile_10_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w60_5 :  std_logic;
signal bh793_w61_5 :  std_logic;
signal bh793_w62_5 :  std_logic;
signal bh793_w63_5 :  std_logic;
signal tile_11_X :  std_logic_vector(3 downto 0);
signal tile_11_Y :  std_logic_vector(0 downto 0);
signal tile_11_output :  std_logic_vector(3 downto 0);
signal tile_11_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w56_5 :  std_logic;
signal bh793_w57_5 :  std_logic;
signal bh793_w58_5 :  std_logic;
signal bh793_w59_5 :  std_logic;
signal tile_12_X :  std_logic_vector(3 downto 0);
signal tile_12_Y :  std_logic_vector(0 downto 0);
signal tile_12_output :  std_logic_vector(3 downto 0);
signal tile_12_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w52_5 :  std_logic;
signal bh793_w53_5 :  std_logic;
signal bh793_w54_5 :  std_logic;
signal bh793_w55_5 :  std_logic;
signal tile_13_X :  std_logic_vector(1 downto 0);
signal tile_13_Y :  std_logic_vector(1 downto 0);
signal tile_13_output :  std_logic_vector(3 downto 0);
signal tile_13_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w65_5 :  std_logic;
signal bh793_w66_5 :  std_logic;
signal bh793_w67_5 :  std_logic;
signal bh793_w68_5 :  std_logic;
signal tile_14_X :  std_logic_vector(2 downto 0);
signal tile_14_Y :  std_logic_vector(1 downto 0);
signal tile_14_output :  std_logic_vector(4 downto 0);
signal tile_14_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w62_6 :  std_logic;
signal bh793_w63_6 :  std_logic;
signal bh793_w64_6 :  std_logic;
signal bh793_w65_6 :  std_logic;
signal bh793_w66_6 :  std_logic;
signal tile_15_X :  std_logic_vector(2 downto 0);
signal tile_15_Y :  std_logic_vector(1 downto 0);
signal tile_15_output :  std_logic_vector(4 downto 0);
signal tile_15_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w59_6 :  std_logic;
signal bh793_w60_6 :  std_logic;
signal bh793_w61_6 :  std_logic;
signal bh793_w62_7 :  std_logic;
signal bh793_w63_7 :  std_logic;
signal tile_16_X :  std_logic_vector(2 downto 0);
signal tile_16_Y :  std_logic_vector(1 downto 0);
signal tile_16_output :  std_logic_vector(4 downto 0);
signal tile_16_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w56_6 :  std_logic;
signal bh793_w57_6 :  std_logic;
signal bh793_w58_6 :  std_logic;
signal bh793_w59_7 :  std_logic;
signal bh793_w60_7 :  std_logic;
signal tile_17_X :  std_logic_vector(2 downto 0);
signal tile_17_Y :  std_logic_vector(1 downto 0);
signal tile_17_output :  std_logic_vector(4 downto 0);
signal tile_17_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w53_6 :  std_logic;
signal bh793_w54_6 :  std_logic;
signal bh793_w55_6 :  std_logic;
signal bh793_w56_7 :  std_logic;
signal bh793_w57_7 :  std_logic;
signal tile_18_X :  std_logic_vector(2 downto 0);
signal tile_18_Y :  std_logic_vector(1 downto 0);
signal tile_18_output :  std_logic_vector(4 downto 0);
signal tile_18_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w50_4 :  std_logic;
signal bh793_w51_5 :  std_logic;
signal bh793_w52_6 :  std_logic;
signal bh793_w53_7 :  std_logic;
signal bh793_w54_7 :  std_logic;
signal tile_19_X :  std_logic_vector(1 downto 0);
signal tile_19_Y :  std_logic_vector(1 downto 0);
signal tile_19_output :  std_logic_vector(3 downto 0);
signal tile_19_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w63_8 :  std_logic;
signal bh793_w64_7 :  std_logic;
signal bh793_w65_7 :  std_logic;
signal bh793_w66_7 :  std_logic;
signal tile_20_X :  std_logic_vector(2 downto 0);
signal tile_20_Y :  std_logic_vector(1 downto 0);
signal tile_20_output :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w60_8 :  std_logic;
signal bh793_w61_7 :  std_logic;
signal bh793_w62_8 :  std_logic;
signal bh793_w63_9 :  std_logic;
signal bh793_w64_8 :  std_logic;
signal tile_21_X :  std_logic_vector(2 downto 0);
signal tile_21_Y :  std_logic_vector(1 downto 0);
signal tile_21_output :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w57_8 :  std_logic;
signal bh793_w58_7 :  std_logic;
signal bh793_w59_8 :  std_logic;
signal bh793_w60_9 :  std_logic;
signal bh793_w61_8 :  std_logic;
signal tile_22_X :  std_logic_vector(2 downto 0);
signal tile_22_Y :  std_logic_vector(1 downto 0);
signal tile_22_output :  std_logic_vector(4 downto 0);
signal tile_22_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w54_8 :  std_logic;
signal bh793_w55_7 :  std_logic;
signal bh793_w56_8 :  std_logic;
signal bh793_w57_9 :  std_logic;
signal bh793_w58_8 :  std_logic;
signal tile_23_X :  std_logic_vector(2 downto 0);
signal tile_23_Y :  std_logic_vector(1 downto 0);
signal tile_23_output :  std_logic_vector(4 downto 0);
signal tile_23_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w51_6 :  std_logic;
signal bh793_w52_7 :  std_logic;
signal bh793_w53_8 :  std_logic;
signal bh793_w54_9 :  std_logic;
signal bh793_w55_8 :  std_logic;
signal tile_24_X :  std_logic_vector(2 downto 0);
signal tile_24_Y :  std_logic_vector(1 downto 0);
signal tile_24_output :  std_logic_vector(4 downto 0);
signal tile_24_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w48_4 :  std_logic;
signal bh793_w49_4 :  std_logic;
signal bh793_w50_5 :  std_logic;
signal bh793_w51_7 :  std_logic;
signal bh793_w52_8 :  std_logic;
signal tile_25_X :  std_logic_vector(0 downto 0);
signal tile_25_Y :  std_logic_vector(0 downto 0);
signal tile_25_output :  std_logic_vector(0 downto 0);
signal tile_25_filtered_output :  std_logic_vector(0 downto 0);
signal bh793_w85_2 :  std_logic;
signal tile_26_X :  std_logic_vector(3 downto 0);
signal tile_26_Y :  std_logic_vector(0 downto 0);
signal tile_26_output :  std_logic_vector(3 downto 0);
signal tile_26_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w81_3 :  std_logic;
signal bh793_w82_2 :  std_logic;
signal bh793_w83_2 :  std_logic;
signal bh793_w84_2 :  std_logic;
signal tile_27_X :  std_logic_vector(3 downto 0);
signal tile_27_Y :  std_logic_vector(0 downto 0);
signal tile_27_output :  std_logic_vector(3 downto 0);
signal tile_27_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w77_3 :  std_logic;
signal bh793_w78_3 :  std_logic;
signal bh793_w79_3 :  std_logic;
signal bh793_w80_3 :  std_logic;
signal tile_28_X :  std_logic_vector(3 downto 0);
signal tile_28_Y :  std_logic_vector(0 downto 0);
signal tile_28_output :  std_logic_vector(3 downto 0);
signal tile_28_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w73_4 :  std_logic;
signal bh793_w74_4 :  std_logic;
signal bh793_w75_4 :  std_logic;
signal bh793_w76_4 :  std_logic;
signal tile_29_X :  std_logic_vector(3 downto 0);
signal tile_29_Y :  std_logic_vector(0 downto 0);
signal tile_29_output :  std_logic_vector(3 downto 0);
signal tile_29_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w69_4 :  std_logic;
signal bh793_w70_4 :  std_logic;
signal bh793_w71_4 :  std_logic;
signal bh793_w72_4 :  std_logic;
signal tile_30_X :  std_logic_vector(1 downto 0);
signal tile_30_Y :  std_logic_vector(1 downto 0);
signal tile_30_output :  std_logic_vector(3 downto 0);
signal tile_30_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w82_3 :  std_logic;
signal bh793_w83_3 :  std_logic;
signal bh793_w84_3 :  std_logic;
signal bh793_w85_3 :  std_logic;
signal tile_31_X :  std_logic_vector(2 downto 0);
signal tile_31_Y :  std_logic_vector(1 downto 0);
signal tile_31_output :  std_logic_vector(4 downto 0);
signal tile_31_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w79_4 :  std_logic;
signal bh793_w80_4 :  std_logic;
signal bh793_w81_4 :  std_logic;
signal bh793_w82_4 :  std_logic;
signal bh793_w83_4 :  std_logic;
signal tile_32_X :  std_logic_vector(2 downto 0);
signal tile_32_Y :  std_logic_vector(1 downto 0);
signal tile_32_output :  std_logic_vector(4 downto 0);
signal tile_32_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w76_5 :  std_logic;
signal bh793_w77_4 :  std_logic;
signal bh793_w78_4 :  std_logic;
signal bh793_w79_5 :  std_logic;
signal bh793_w80_5 :  std_logic;
signal tile_33_X :  std_logic_vector(2 downto 0);
signal tile_33_Y :  std_logic_vector(1 downto 0);
signal tile_33_output :  std_logic_vector(4 downto 0);
signal tile_33_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w73_5 :  std_logic;
signal bh793_w74_5 :  std_logic;
signal bh793_w75_5 :  std_logic;
signal bh793_w76_6 :  std_logic;
signal bh793_w77_5 :  std_logic;
signal tile_34_X :  std_logic_vector(2 downto 0);
signal tile_34_Y :  std_logic_vector(1 downto 0);
signal tile_34_output :  std_logic_vector(4 downto 0);
signal tile_34_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w70_5 :  std_logic;
signal bh793_w71_5 :  std_logic;
signal bh793_w72_5 :  std_logic;
signal bh793_w73_6 :  std_logic;
signal bh793_w74_6 :  std_logic;
signal tile_35_X :  std_logic_vector(2 downto 0);
signal tile_35_Y :  std_logic_vector(1 downto 0);
signal tile_35_output :  std_logic_vector(4 downto 0);
signal tile_35_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w67_6 :  std_logic;
signal bh793_w68_6 :  std_logic;
signal bh793_w69_5 :  std_logic;
signal bh793_w70_6 :  std_logic;
signal bh793_w71_6 :  std_logic;
signal tile_36_X :  std_logic_vector(1 downto 0);
signal tile_36_Y :  std_logic_vector(1 downto 0);
signal tile_36_output :  std_logic_vector(3 downto 0);
signal tile_36_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w80_6 :  std_logic;
signal bh793_w81_5 :  std_logic;
signal bh793_w82_5 :  std_logic;
signal bh793_w83_5 :  std_logic;
signal tile_37_X :  std_logic_vector(2 downto 0);
signal tile_37_Y :  std_logic_vector(1 downto 0);
signal tile_37_output :  std_logic_vector(4 downto 0);
signal tile_37_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w77_6 :  std_logic;
signal bh793_w78_5 :  std_logic;
signal bh793_w79_6 :  std_logic;
signal bh793_w80_7 :  std_logic;
signal bh793_w81_6 :  std_logic;
signal tile_38_X :  std_logic_vector(2 downto 0);
signal tile_38_Y :  std_logic_vector(1 downto 0);
signal tile_38_output :  std_logic_vector(4 downto 0);
signal tile_38_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w74_7 :  std_logic;
signal bh793_w75_6 :  std_logic;
signal bh793_w76_7 :  std_logic;
signal bh793_w77_7 :  std_logic;
signal bh793_w78_6 :  std_logic;
signal tile_39_X :  std_logic_vector(2 downto 0);
signal tile_39_Y :  std_logic_vector(1 downto 0);
signal tile_39_output :  std_logic_vector(4 downto 0);
signal tile_39_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w71_7 :  std_logic;
signal bh793_w72_6 :  std_logic;
signal bh793_w73_7 :  std_logic;
signal bh793_w74_8 :  std_logic;
signal bh793_w75_7 :  std_logic;
signal tile_40_X :  std_logic_vector(2 downto 0);
signal tile_40_Y :  std_logic_vector(1 downto 0);
signal tile_40_output :  std_logic_vector(4 downto 0);
signal tile_40_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w68_7 :  std_logic;
signal bh793_w69_6 :  std_logic;
signal bh793_w70_7 :  std_logic;
signal bh793_w71_8 :  std_logic;
signal bh793_w72_7 :  std_logic;
signal tile_41_X :  std_logic_vector(2 downto 0);
signal tile_41_Y :  std_logic_vector(1 downto 0);
signal tile_41_output :  std_logic_vector(4 downto 0);
signal tile_41_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w65_8 :  std_logic;
signal bh793_w66_8 :  std_logic;
signal bh793_w67_7 :  std_logic;
signal bh793_w68_8 :  std_logic;
signal bh793_w69_7 :  std_logic;
signal tile_42_X :  std_logic_vector(0 downto 0);
signal tile_42_Y :  std_logic_vector(0 downto 0);
signal tile_42_output :  std_logic_vector(0 downto 0);
signal tile_42_filtered_output :  std_logic_vector(0 downto 0);
signal bh793_w102_0 :  std_logic;
signal tile_43_X :  std_logic_vector(3 downto 0);
signal tile_43_Y :  std_logic_vector(0 downto 0);
signal tile_43_output :  std_logic_vector(3 downto 0);
signal tile_43_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w98_2 :  std_logic;
signal bh793_w99_1 :  std_logic;
signal bh793_w100_1 :  std_logic;
signal bh793_w101_0 :  std_logic;
signal tile_44_X :  std_logic_vector(3 downto 0);
signal tile_44_Y :  std_logic_vector(0 downto 0);
signal tile_44_output :  std_logic_vector(3 downto 0);
signal tile_44_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w94_2 :  std_logic;
signal bh793_w95_2 :  std_logic;
signal bh793_w96_2 :  std_logic;
signal bh793_w97_2 :  std_logic;
signal tile_45_X :  std_logic_vector(3 downto 0);
signal tile_45_Y :  std_logic_vector(0 downto 0);
signal tile_45_output :  std_logic_vector(3 downto 0);
signal tile_45_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w90_2 :  std_logic;
signal bh793_w91_2 :  std_logic;
signal bh793_w92_2 :  std_logic;
signal bh793_w93_2 :  std_logic;
signal tile_46_X :  std_logic_vector(3 downto 0);
signal tile_46_Y :  std_logic_vector(0 downto 0);
signal tile_46_output :  std_logic_vector(3 downto 0);
signal tile_46_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w86_2 :  std_logic;
signal bh793_w87_2 :  std_logic;
signal bh793_w88_2 :  std_logic;
signal bh793_w89_2 :  std_logic;
signal tile_47_X :  std_logic_vector(1 downto 0);
signal tile_47_Y :  std_logic_vector(1 downto 0);
signal tile_47_output :  std_logic_vector(3 downto 0);
signal tile_47_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w99_2 :  std_logic;
signal bh793_w100_2 :  std_logic;
signal bh793_w101_1 :  std_logic;
signal bh793_w102_1 :  std_logic;
signal tile_48_X :  std_logic_vector(2 downto 0);
signal tile_48_Y :  std_logic_vector(1 downto 0);
signal tile_48_output :  std_logic_vector(4 downto 0);
signal tile_48_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w96_3 :  std_logic;
signal bh793_w97_3 :  std_logic;
signal bh793_w98_3 :  std_logic;
signal bh793_w99_3 :  std_logic;
signal bh793_w100_3 :  std_logic;
signal tile_49_X :  std_logic_vector(2 downto 0);
signal tile_49_Y :  std_logic_vector(1 downto 0);
signal tile_49_output :  std_logic_vector(4 downto 0);
signal tile_49_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w93_3 :  std_logic;
signal bh793_w94_3 :  std_logic;
signal bh793_w95_3 :  std_logic;
signal bh793_w96_4 :  std_logic;
signal bh793_w97_4 :  std_logic;
signal tile_50_X :  std_logic_vector(2 downto 0);
signal tile_50_Y :  std_logic_vector(1 downto 0);
signal tile_50_output :  std_logic_vector(4 downto 0);
signal tile_50_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w90_3 :  std_logic;
signal bh793_w91_3 :  std_logic;
signal bh793_w92_3 :  std_logic;
signal bh793_w93_4 :  std_logic;
signal bh793_w94_4 :  std_logic;
signal tile_51_X :  std_logic_vector(2 downto 0);
signal tile_51_Y :  std_logic_vector(1 downto 0);
signal tile_51_output :  std_logic_vector(4 downto 0);
signal tile_51_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w87_3 :  std_logic;
signal bh793_w88_3 :  std_logic;
signal bh793_w89_3 :  std_logic;
signal bh793_w90_4 :  std_logic;
signal bh793_w91_4 :  std_logic;
signal tile_52_X :  std_logic_vector(2 downto 0);
signal tile_52_Y :  std_logic_vector(1 downto 0);
signal tile_52_output :  std_logic_vector(4 downto 0);
signal tile_52_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w84_4 :  std_logic;
signal bh793_w85_4 :  std_logic;
signal bh793_w86_3 :  std_logic;
signal bh793_w87_4 :  std_logic;
signal bh793_w88_4 :  std_logic;
signal tile_53_X :  std_logic_vector(1 downto 0);
signal tile_53_Y :  std_logic_vector(1 downto 0);
signal tile_53_output :  std_logic_vector(3 downto 0);
signal tile_53_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w97_5 :  std_logic;
signal bh793_w98_4 :  std_logic;
signal bh793_w99_4 :  std_logic;
signal bh793_w100_4 :  std_logic;
signal tile_54_X :  std_logic_vector(2 downto 0);
signal tile_54_Y :  std_logic_vector(1 downto 0);
signal tile_54_output :  std_logic_vector(4 downto 0);
signal tile_54_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w94_5 :  std_logic;
signal bh793_w95_4 :  std_logic;
signal bh793_w96_5 :  std_logic;
signal bh793_w97_6 :  std_logic;
signal bh793_w98_5 :  std_logic;
signal tile_55_X :  std_logic_vector(2 downto 0);
signal tile_55_Y :  std_logic_vector(1 downto 0);
signal tile_55_output :  std_logic_vector(4 downto 0);
signal tile_55_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w91_5 :  std_logic;
signal bh793_w92_4 :  std_logic;
signal bh793_w93_5 :  std_logic;
signal bh793_w94_6 :  std_logic;
signal bh793_w95_5 :  std_logic;
signal tile_56_X :  std_logic_vector(2 downto 0);
signal tile_56_Y :  std_logic_vector(1 downto 0);
signal tile_56_output :  std_logic_vector(4 downto 0);
signal tile_56_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w88_5 :  std_logic;
signal bh793_w89_4 :  std_logic;
signal bh793_w90_5 :  std_logic;
signal bh793_w91_6 :  std_logic;
signal bh793_w92_5 :  std_logic;
signal tile_57_X :  std_logic_vector(2 downto 0);
signal tile_57_Y :  std_logic_vector(1 downto 0);
signal tile_57_output :  std_logic_vector(4 downto 0);
signal tile_57_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w85_5 :  std_logic;
signal bh793_w86_4 :  std_logic;
signal bh793_w87_5 :  std_logic;
signal bh793_w88_6 :  std_logic;
signal bh793_w89_5 :  std_logic;
signal tile_58_X :  std_logic_vector(2 downto 0);
signal tile_58_Y :  std_logic_vector(1 downto 0);
signal tile_58_output :  std_logic_vector(4 downto 0);
signal tile_58_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w82_6 :  std_logic;
signal bh793_w83_6 :  std_logic;
signal bh793_w84_5 :  std_logic;
signal bh793_w85_6 :  std_logic;
signal bh793_w86_5 :  std_logic;
signal tile_59_X :  std_logic_vector(1 downto 0);
signal tile_59_Y :  std_logic_vector(1 downto 0);
signal tile_59_output :  std_logic_vector(3 downto 0);
signal tile_59_filtered_output :  std_logic_vector(3 downto 0);
signal bh793_w102_2 :  std_logic;
signal bh793_w103_0 :  std_logic;
signal bh793_w104_0 :  std_logic;
signal bh793_w105_0 :  std_logic;
signal tile_60_X :  std_logic_vector(1 downto 0);
signal tile_60_Y :  std_logic_vector(2 downto 0);
signal tile_60_output :  std_logic_vector(4 downto 0);
signal tile_60_filtered_output :  std_logic_vector(4 downto 0);
signal bh793_w99_5 :  std_logic;
signal bh793_w100_5 :  std_logic;
signal bh793_w101_2 :  std_logic;
signal bh793_w102_3 :  std_logic;
signal bh793_w103_1 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1033_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1033_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1033_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1033_Out0_copy1034 :  std_logic_vector(2 downto 0);
signal bh793_w17_2 :  std_logic;
signal bh793_w18_2 :  std_logic;
signal bh793_w19_2 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1035_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1035_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1035_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1035_Out0_copy1036 :  std_logic_vector(2 downto 0);
signal bh793_w19_3 :  std_logic;
signal bh793_w20_2 :  std_logic;
signal bh793_w21_2 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1037_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1037_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1037_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1037_Out0_copy1038 :  std_logic_vector(2 downto 0);
signal bh793_w21_3 :  std_logic;
signal bh793_w22_2 :  std_logic;
signal bh793_w23_2 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1041_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1041_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1041_Out0_copy1042 :  std_logic_vector(1 downto 0);
signal bh793_w23_3 :  std_logic;
signal bh793_w24_3 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1043_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1043_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1043_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1043_Out0_copy1044 :  std_logic_vector(2 downto 0);
signal bh793_w24_4 :  std_logic;
signal bh793_w25_3 :  std_logic;
signal bh793_w26_3 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1045_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1045_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1045_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1045_Out0_copy1046 :  std_logic_vector(2 downto 0);
signal bh793_w26_4 :  std_logic;
signal bh793_w27_3 :  std_logic;
signal bh793_w28_3 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1047_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1047_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1047_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1047_Out0_copy1048 :  std_logic_vector(2 downto 0);
signal bh793_w28_4 :  std_logic;
signal bh793_w29_3 :  std_logic;
signal bh793_w30_3 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1049_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1049_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1049_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1049_Out0_copy1050 :  std_logic_vector(2 downto 0);
signal bh793_w30_4 :  std_logic;
signal bh793_w31_3 :  std_logic;
signal bh793_w32_3 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1051_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1051_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1051_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1051_Out0_copy1052 :  std_logic_vector(2 downto 0);
signal bh793_w32_4 :  std_logic;
signal bh793_w33_3 :  std_logic;
signal bh793_w34_4 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1055_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1055_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1055_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1055_Out0_copy1056 :  std_logic_vector(2 downto 0);
signal bh793_w34_5 :  std_logic;
signal bh793_w35_4 :  std_logic;
signal bh793_w36_4 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1057_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1057_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1057_Out0_copy1058 :  std_logic_vector(1 downto 0);
signal bh793_w35_5 :  std_logic;
signal bh793_w36_5 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1059_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1059_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1059_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1059_Out0_copy1060 :  std_logic_vector(2 downto 0);
signal bh793_w36_6 :  std_logic;
signal bh793_w37_4 :  std_logic;
signal bh793_w38_4 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1061_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1061_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1061_Out0_copy1062 :  std_logic_vector(1 downto 0);
signal bh793_w37_5 :  std_logic;
signal bh793_w38_5 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1063_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1063_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1063_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1063_Out0_copy1064 :  std_logic_vector(2 downto 0);
signal bh793_w38_6 :  std_logic;
signal bh793_w39_4 :  std_logic;
signal bh793_w40_4 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1065_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1065_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1065_Out0_copy1066 :  std_logic_vector(1 downto 0);
signal bh793_w39_5 :  std_logic;
signal bh793_w40_5 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1067_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1067_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1067_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1067_Out0_copy1068 :  std_logic_vector(2 downto 0);
signal bh793_w40_6 :  std_logic;
signal bh793_w41_4 :  std_logic;
signal bh793_w42_4 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1069_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1069_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1069_Out0_copy1070 :  std_logic_vector(1 downto 0);
signal bh793_w41_5 :  std_logic;
signal bh793_w42_5 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1071_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1071_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1071_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1071_Out0_copy1072 :  std_logic_vector(2 downto 0);
signal bh793_w42_6 :  std_logic;
signal bh793_w43_4 :  std_logic;
signal bh793_w44_4 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1073_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1073_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1073_Out0_copy1074 :  std_logic_vector(1 downto 0);
signal bh793_w43_5 :  std_logic;
signal bh793_w44_5 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1075_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1075_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1075_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1075_Out0_copy1076 :  std_logic_vector(2 downto 0);
signal bh793_w44_6 :  std_logic;
signal bh793_w45_4 :  std_logic;
signal bh793_w46_4 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1077_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1077_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1077_Out0_copy1078 :  std_logic_vector(1 downto 0);
signal bh793_w45_5 :  std_logic;
signal bh793_w46_5 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1079_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1079_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1079_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1079_Out0_copy1080 :  std_logic_vector(2 downto 0);
signal bh793_w46_6 :  std_logic;
signal bh793_w47_4 :  std_logic;
signal bh793_w48_5 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1081_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1081_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1081_Out0_copy1082 :  std_logic_vector(1 downto 0);
signal bh793_w47_5 :  std_logic;
signal bh793_w48_6 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1083_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1083_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1083_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1083_Out0_copy1084 :  std_logic_vector(2 downto 0);
signal bh793_w48_7 :  std_logic;
signal bh793_w49_5 :  std_logic;
signal bh793_w50_6 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1085_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1085_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1085_Out0_copy1086 :  std_logic_vector(1 downto 0);
signal bh793_w49_6 :  std_logic;
signal bh793_w50_7 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1089_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1089_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1089_Out0_copy1090 :  std_logic_vector(2 downto 0);
signal bh793_w50_8 :  std_logic;
signal bh793_w51_8 :  std_logic;
signal bh793_w52_9 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1091_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1091_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1091_Out0_copy1092 :  std_logic_vector(2 downto 0);
signal bh793_w51_9 :  std_logic;
signal bh793_w52_10 :  std_logic;
signal bh793_w53_9 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1093_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1093_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1093_Out0_copy1094 :  std_logic_vector(1 downto 0);
signal bh793_w51_10 :  std_logic;
signal bh793_w52_11 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1095_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1095_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1095_Out0_copy1096 :  std_logic_vector(2 downto 0);
signal bh793_w52_12 :  std_logic;
signal bh793_w53_10 :  std_logic;
signal bh793_w54_10 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1097_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1097_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1097_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1097_Out0_copy1098 :  std_logic_vector(2 downto 0);
signal bh793_w52_13 :  std_logic;
signal bh793_w53_11 :  std_logic;
signal bh793_w54_11 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1099_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1099_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1099_Out0_copy1100 :  std_logic_vector(2 downto 0);
signal bh793_w53_12 :  std_logic;
signal bh793_w54_12 :  std_logic;
signal bh793_w55_9 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1101_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1101_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1101_Out0_copy1102 :  std_logic_vector(2 downto 0);
signal bh793_w54_13 :  std_logic;
signal bh793_w55_10 :  std_logic;
signal bh793_w56_9 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1103_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1103_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1103_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1103_Out0_copy1104 :  std_logic_vector(2 downto 0);
signal bh793_w54_14 :  std_logic;
signal bh793_w55_11 :  std_logic;
signal bh793_w56_10 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1105_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1105_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1105_Out0_copy1106 :  std_logic_vector(2 downto 0);
signal bh793_w55_12 :  std_logic;
signal bh793_w56_11 :  std_logic;
signal bh793_w57_10 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1107_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1107_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1107_Out0_copy1108 :  std_logic_vector(1 downto 0);
signal bh793_w55_13 :  std_logic;
signal bh793_w56_12 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1109_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1109_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1109_Out0_copy1110 :  std_logic_vector(2 downto 0);
signal bh793_w56_13 :  std_logic;
signal bh793_w57_11 :  std_logic;
signal bh793_w58_9 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1111_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1111_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1111_Out0_copy1112 :  std_logic_vector(1 downto 0);
signal bh793_w56_14 :  std_logic;
signal bh793_w57_12 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1113_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1113_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1113_Out0_copy1114 :  std_logic_vector(2 downto 0);
signal bh793_w57_13 :  std_logic;
signal bh793_w58_10 :  std_logic;
signal bh793_w59_9 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1115_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1115_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1115_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1115_Out0_copy1116 :  std_logic_vector(2 downto 0);
signal bh793_w57_14 :  std_logic;
signal bh793_w58_11 :  std_logic;
signal bh793_w59_10 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1117_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1117_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1117_Out0_copy1118 :  std_logic_vector(2 downto 0);
signal bh793_w58_12 :  std_logic;
signal bh793_w59_11 :  std_logic;
signal bh793_w60_10 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1119_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1119_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1119_Out0_copy1120 :  std_logic_vector(1 downto 0);
signal bh793_w58_13 :  std_logic;
signal bh793_w59_12 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1121_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1121_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1121_Out0_copy1122 :  std_logic_vector(2 downto 0);
signal bh793_w59_13 :  std_logic;
signal bh793_w60_11 :  std_logic;
signal bh793_w61_9 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1123_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1123_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1123_Out0_copy1124 :  std_logic_vector(1 downto 0);
signal bh793_w59_14 :  std_logic;
signal bh793_w60_12 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1125_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1125_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1125_Out0_copy1126 :  std_logic_vector(2 downto 0);
signal bh793_w60_13 :  std_logic;
signal bh793_w61_10 :  std_logic;
signal bh793_w62_9 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1127_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1127_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1127_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1127_Out0_copy1128 :  std_logic_vector(2 downto 0);
signal bh793_w60_14 :  std_logic;
signal bh793_w61_11 :  std_logic;
signal bh793_w62_10 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1129_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1129_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1129_Out0_copy1130 :  std_logic_vector(2 downto 0);
signal bh793_w61_12 :  std_logic;
signal bh793_w62_11 :  std_logic;
signal bh793_w63_10 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1131_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1131_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1131_Out0_copy1132 :  std_logic_vector(1 downto 0);
signal bh793_w61_13 :  std_logic;
signal bh793_w62_12 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1133_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1133_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1133_Out0_copy1134 :  std_logic_vector(2 downto 0);
signal bh793_w62_13 :  std_logic;
signal bh793_w63_11 :  std_logic;
signal bh793_w64_9 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1135_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1135_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1135_Out0_copy1136 :  std_logic_vector(1 downto 0);
signal bh793_w62_14 :  std_logic;
signal bh793_w63_12 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1137_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1137_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1137_Out0_copy1138 :  std_logic_vector(2 downto 0);
signal bh793_w63_13 :  std_logic;
signal bh793_w64_10 :  std_logic;
signal bh793_w65_9 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1139_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1139_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1139_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1139_Out0_copy1140 :  std_logic_vector(2 downto 0);
signal bh793_w63_14 :  std_logic;
signal bh793_w64_11 :  std_logic;
signal bh793_w65_10 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1141_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1141_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1141_Out0_copy1142 :  std_logic_vector(2 downto 0);
signal bh793_w64_12 :  std_logic;
signal bh793_w65_11 :  std_logic;
signal bh793_w66_9 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1143_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1143_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1143_Out0_copy1144 :  std_logic_vector(1 downto 0);
signal bh793_w64_13 :  std_logic;
signal bh793_w65_12 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1145_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1145_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1145_Out0_copy1146 :  std_logic_vector(2 downto 0);
signal bh793_w65_13 :  std_logic;
signal bh793_w66_10 :  std_logic;
signal bh793_w67_8 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1147_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1147_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1147_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1147_Out0_copy1148 :  std_logic_vector(2 downto 0);
signal bh793_w65_14 :  std_logic;
signal bh793_w66_11 :  std_logic;
signal bh793_w67_9 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1149_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1149_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1149_Out0_copy1150 :  std_logic_vector(2 downto 0);
signal bh793_w66_12 :  std_logic;
signal bh793_w67_10 :  std_logic;
signal bh793_w68_9 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1151_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1151_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1151_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1151_Out0_copy1152 :  std_logic_vector(2 downto 0);
signal bh793_w66_13 :  std_logic;
signal bh793_w67_11 :  std_logic;
signal bh793_w68_10 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1153_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1153_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1153_Out0_copy1154 :  std_logic_vector(2 downto 0);
signal bh793_w67_12 :  std_logic;
signal bh793_w68_11 :  std_logic;
signal bh793_w69_8 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1155_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1155_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1155_Out0_copy1156 :  std_logic_vector(2 downto 0);
signal bh793_w68_12 :  std_logic;
signal bh793_w69_9 :  std_logic;
signal bh793_w70_8 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1157_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1157_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1157_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1157_Out0_copy1158 :  std_logic_vector(2 downto 0);
signal bh793_w68_13 :  std_logic;
signal bh793_w69_10 :  std_logic;
signal bh793_w70_9 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1159_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1159_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1159_Out0_copy1160 :  std_logic_vector(2 downto 0);
signal bh793_w69_11 :  std_logic;
signal bh793_w70_10 :  std_logic;
signal bh793_w71_9 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1161_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1161_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1161_Out0_copy1162 :  std_logic_vector(2 downto 0);
signal bh793_w70_11 :  std_logic;
signal bh793_w71_10 :  std_logic;
signal bh793_w72_8 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1163_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1163_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1163_Out0_copy1164 :  std_logic_vector(1 downto 0);
signal bh793_w70_12 :  std_logic;
signal bh793_w71_11 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1165_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1165_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1165_Out0_copy1166 :  std_logic_vector(2 downto 0);
signal bh793_w71_12 :  std_logic;
signal bh793_w72_9 :  std_logic;
signal bh793_w73_8 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1167_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1167_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1167_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1167_Out0_copy1168 :  std_logic_vector(2 downto 0);
signal bh793_w71_13 :  std_logic;
signal bh793_w72_10 :  std_logic;
signal bh793_w73_9 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1169_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1169_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1169_Out0_copy1170 :  std_logic_vector(2 downto 0);
signal bh793_w72_11 :  std_logic;
signal bh793_w73_10 :  std_logic;
signal bh793_w74_9 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1171_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1171_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1171_Out0_copy1172 :  std_logic_vector(2 downto 0);
signal bh793_w73_11 :  std_logic;
signal bh793_w74_10 :  std_logic;
signal bh793_w75_8 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1173_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1173_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1173_Out0_copy1174 :  std_logic_vector(1 downto 0);
signal bh793_w73_12 :  std_logic;
signal bh793_w74_11 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1175_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1175_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1175_Out0_copy1176 :  std_logic_vector(2 downto 0);
signal bh793_w74_12 :  std_logic;
signal bh793_w75_9 :  std_logic;
signal bh793_w76_8 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1177_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1177_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1177_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1177_Out0_copy1178 :  std_logic_vector(2 downto 0);
signal bh793_w74_13 :  std_logic;
signal bh793_w75_10 :  std_logic;
signal bh793_w76_9 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1179_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1179_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1179_Out0_copy1180 :  std_logic_vector(2 downto 0);
signal bh793_w75_11 :  std_logic;
signal bh793_w76_10 :  std_logic;
signal bh793_w77_8 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1181_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1181_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1181_Out0_copy1182 :  std_logic_vector(2 downto 0);
signal bh793_w76_11 :  std_logic;
signal bh793_w77_9 :  std_logic;
signal bh793_w78_7 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1183_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1183_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1183_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1183_Out0_copy1184 :  std_logic_vector(2 downto 0);
signal bh793_w76_12 :  std_logic;
signal bh793_w77_10 :  std_logic;
signal bh793_w78_8 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1185_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1185_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1185_Out0_copy1186 :  std_logic_vector(2 downto 0);
signal bh793_w77_11 :  std_logic;
signal bh793_w78_9 :  std_logic;
signal bh793_w79_7 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1187_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1187_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1187_Out0_copy1188 :  std_logic_vector(2 downto 0);
signal bh793_w78_10 :  std_logic;
signal bh793_w79_8 :  std_logic;
signal bh793_w80_8 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1189_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1189_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1189_Out0_copy1190 :  std_logic_vector(2 downto 0);
signal bh793_w79_9 :  std_logic;
signal bh793_w80_9 :  std_logic;
signal bh793_w81_7 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1191_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1191_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1191_Out0_copy1192 :  std_logic_vector(2 downto 0);
signal bh793_w80_10 :  std_logic;
signal bh793_w81_8 :  std_logic;
signal bh793_w82_7 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1193_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1193_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1193_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1193_Out0_copy1194 :  std_logic_vector(2 downto 0);
signal bh793_w80_11 :  std_logic;
signal bh793_w81_9 :  std_logic;
signal bh793_w82_8 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1195_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1195_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1195_Out0_copy1196 :  std_logic_vector(2 downto 0);
signal bh793_w81_10 :  std_logic;
signal bh793_w82_9 :  std_logic;
signal bh793_w83_7 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1197_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1197_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1197_Out0_copy1198 :  std_logic_vector(2 downto 0);
signal bh793_w82_10 :  std_logic;
signal bh793_w83_8 :  std_logic;
signal bh793_w84_6 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1199_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1199_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1199_Out0_copy1200 :  std_logic_vector(2 downto 0);
signal bh793_w83_9 :  std_logic;
signal bh793_w84_7 :  std_logic;
signal bh793_w85_7 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1201_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1201_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1201_Out0_copy1202 :  std_logic_vector(2 downto 0);
signal bh793_w84_8 :  std_logic;
signal bh793_w85_8 :  std_logic;
signal bh793_w86_6 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1203_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1203_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1203_Out0_copy1204 :  std_logic_vector(2 downto 0);
signal bh793_w85_9 :  std_logic;
signal bh793_w86_7 :  std_logic;
signal bh793_w87_6 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1205_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1205_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1205_Out0_copy1206 :  std_logic_vector(2 downto 0);
signal bh793_w86_8 :  std_logic;
signal bh793_w87_7 :  std_logic;
signal bh793_w88_7 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1207_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1207_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1207_Out0_copy1208 :  std_logic_vector(2 downto 0);
signal bh793_w87_8 :  std_logic;
signal bh793_w88_8 :  std_logic;
signal bh793_w89_6 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1209_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1209_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1209_Out0_copy1210 :  std_logic_vector(2 downto 0);
signal bh793_w88_9 :  std_logic;
signal bh793_w89_7 :  std_logic;
signal bh793_w90_6 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1211_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1211_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1211_Out0_copy1212 :  std_logic_vector(2 downto 0);
signal bh793_w89_8 :  std_logic;
signal bh793_w90_7 :  std_logic;
signal bh793_w91_7 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1213_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1213_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1213_Out0_copy1214 :  std_logic_vector(2 downto 0);
signal bh793_w90_8 :  std_logic;
signal bh793_w91_8 :  std_logic;
signal bh793_w92_6 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1215_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1215_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1215_Out0_copy1216 :  std_logic_vector(2 downto 0);
signal bh793_w91_9 :  std_logic;
signal bh793_w92_7 :  std_logic;
signal bh793_w93_6 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1217_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1217_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1217_Out0_copy1218 :  std_logic_vector(2 downto 0);
signal bh793_w92_8 :  std_logic;
signal bh793_w93_7 :  std_logic;
signal bh793_w94_7 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1219_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1219_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1219_Out0_copy1220 :  std_logic_vector(2 downto 0);
signal bh793_w93_8 :  std_logic;
signal bh793_w94_8 :  std_logic;
signal bh793_w95_6 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1221_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1221_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1221_Out0_copy1222 :  std_logic_vector(2 downto 0);
signal bh793_w94_9 :  std_logic;
signal bh793_w95_7 :  std_logic;
signal bh793_w96_6 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1223_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1223_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1223_Out0_copy1224 :  std_logic_vector(2 downto 0);
signal bh793_w95_8 :  std_logic;
signal bh793_w96_7 :  std_logic;
signal bh793_w97_7 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1225_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1225_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1225_Out0_copy1226 :  std_logic_vector(2 downto 0);
signal bh793_w96_8 :  std_logic;
signal bh793_w97_8 :  std_logic;
signal bh793_w98_6 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1227_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1227_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1227_Out0_copy1228 :  std_logic_vector(2 downto 0);
signal bh793_w97_9 :  std_logic;
signal bh793_w98_7 :  std_logic;
signal bh793_w99_6 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1229_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1229_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1229_Out0_copy1230 :  std_logic_vector(2 downto 0);
signal bh793_w98_8 :  std_logic;
signal bh793_w99_7 :  std_logic;
signal bh793_w100_6 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1231_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1231_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1231_Out0_copy1232 :  std_logic_vector(2 downto 0);
signal bh793_w99_8 :  std_logic;
signal bh793_w100_7 :  std_logic;
signal bh793_w101_3 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1233_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1233_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1233_Out0_copy1234 :  std_logic_vector(2 downto 0);
signal bh793_w100_8 :  std_logic;
signal bh793_w101_4 :  std_logic;
signal bh793_w102_4 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1235_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1235_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1235_Out0_copy1236 :  std_logic_vector(1 downto 0);
signal bh793_w101_5 :  std_logic;
signal bh793_w102_5 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1237_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1237_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1237_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1237_Out0_copy1238 :  std_logic_vector(2 downto 0);
signal bh793_w102_6 :  std_logic;
signal bh793_w103_2 :  std_logic;
signal bh793_w104_1 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1239_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1239_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1239_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1239_Out0_copy1240 :  std_logic_vector(2 downto 0);
signal bh793_w19_4 :  std_logic;
signal bh793_w20_3 :  std_logic;
signal bh793_w21_4 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1241_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1241_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1241_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1241_Out0_copy1242 :  std_logic_vector(2 downto 0);
signal bh793_w21_5 :  std_logic;
signal bh793_w22_3 :  std_logic;
signal bh793_w23_4 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1243_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1243_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1243_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1243_Out0_copy1244 :  std_logic_vector(2 downto 0);
signal bh793_w23_5 :  std_logic;
signal bh793_w24_5 :  std_logic;
signal bh793_w25_4 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1245_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1245_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1245_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1245_Out0_copy1246 :  std_logic_vector(2 downto 0);
signal bh793_w25_5 :  std_logic;
signal bh793_w26_5 :  std_logic;
signal bh793_w27_4 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1247_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1247_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1247_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1247_Out0_copy1248 :  std_logic_vector(2 downto 0);
signal bh793_w27_5 :  std_logic;
signal bh793_w28_5 :  std_logic;
signal bh793_w29_4 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1249_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1249_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1249_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1249_Out0_copy1250 :  std_logic_vector(2 downto 0);
signal bh793_w29_5 :  std_logic;
signal bh793_w30_5 :  std_logic;
signal bh793_w31_4 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1251_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1251_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1251_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1251_Out0_copy1252 :  std_logic_vector(2 downto 0);
signal bh793_w31_5 :  std_logic;
signal bh793_w32_5 :  std_logic;
signal bh793_w33_4 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1253_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1253_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1253_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1253_Out0_copy1254 :  std_logic_vector(2 downto 0);
signal bh793_w33_5 :  std_logic;
signal bh793_w34_6 :  std_logic;
signal bh793_w35_6 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1255_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1255_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1255_Out0_copy1256 :  std_logic_vector(1 downto 0);
signal bh793_w35_7 :  std_logic;
signal bh793_w36_7 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1257_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1257_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1257_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1257_Out0_copy1258 :  std_logic_vector(2 downto 0);
signal bh793_w36_8 :  std_logic;
signal bh793_w37_6 :  std_logic;
signal bh793_w38_7 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1259_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1259_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1259_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1259_Out0_copy1260 :  std_logic_vector(2 downto 0);
signal bh793_w38_8 :  std_logic;
signal bh793_w39_6 :  std_logic;
signal bh793_w40_7 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1261_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1261_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1261_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1261_Out0_copy1262 :  std_logic_vector(2 downto 0);
signal bh793_w40_8 :  std_logic;
signal bh793_w41_6 :  std_logic;
signal bh793_w42_7 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1263_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1263_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1263_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1263_Out0_copy1264 :  std_logic_vector(2 downto 0);
signal bh793_w42_8 :  std_logic;
signal bh793_w43_6 :  std_logic;
signal bh793_w44_7 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1265_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1265_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1265_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1265_Out0_copy1266 :  std_logic_vector(2 downto 0);
signal bh793_w44_8 :  std_logic;
signal bh793_w45_6 :  std_logic;
signal bh793_w46_7 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1267_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1267_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1267_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1267_Out0_copy1268 :  std_logic_vector(2 downto 0);
signal bh793_w46_8 :  std_logic;
signal bh793_w47_6 :  std_logic;
signal bh793_w48_8 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1269_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1269_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1269_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1269_Out0_copy1270 :  std_logic_vector(2 downto 0);
signal bh793_w48_9 :  std_logic;
signal bh793_w49_7 :  std_logic;
signal bh793_w50_9 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1271_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1271_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1271_Out0_copy1272 :  std_logic_vector(1 downto 0);
signal bh793_w49_8 :  std_logic;
signal bh793_w50_10 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1273_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1273_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1273_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1273_Out0_copy1274 :  std_logic_vector(2 downto 0);
signal bh793_w50_11 :  std_logic;
signal bh793_w51_11 :  std_logic;
signal bh793_w52_14 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1275_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1275_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1275_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1275_Out0_copy1276 :  std_logic_vector(2 downto 0);
signal bh793_w52_15 :  std_logic;
signal bh793_w53_13 :  std_logic;
signal bh793_w54_15 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1277_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1277_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1277_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1277_Out0_copy1278 :  std_logic_vector(2 downto 0);
signal bh793_w53_14 :  std_logic;
signal bh793_w54_16 :  std_logic;
signal bh793_w55_14 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1279_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1279_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1279_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1279_Out0_copy1280 :  std_logic_vector(2 downto 0);
signal bh793_w54_17 :  std_logic;
signal bh793_w55_15 :  std_logic;
signal bh793_w56_15 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1281_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1281_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1281_Out0_copy1282 :  std_logic_vector(1 downto 0);
signal bh793_w55_16 :  std_logic;
signal bh793_w56_16 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1283_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1283_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1283_Out0_copy1284 :  std_logic_vector(2 downto 0);
signal bh793_w56_17 :  std_logic;
signal bh793_w57_15 :  std_logic;
signal bh793_w58_14 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1285_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1285_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1285_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1285_Out0_copy1286 :  std_logic_vector(2 downto 0);
signal bh793_w57_16 :  std_logic;
signal bh793_w58_15 :  std_logic;
signal bh793_w59_15 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1287_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1287_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1287_Out0_copy1288 :  std_logic_vector(1 downto 0);
signal bh793_w58_16 :  std_logic;
signal bh793_w59_16 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1289_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1289_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1289_Out0_copy1290 :  std_logic_vector(2 downto 0);
signal bh793_w59_17 :  std_logic;
signal bh793_w60_15 :  std_logic;
signal bh793_w61_14 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1291_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1291_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1291_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1291_Out0_copy1292 :  std_logic_vector(2 downto 0);
signal bh793_w60_16 :  std_logic;
signal bh793_w61_15 :  std_logic;
signal bh793_w62_15 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1293_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1293_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1293_Out0_copy1294 :  std_logic_vector(1 downto 0);
signal bh793_w61_16 :  std_logic;
signal bh793_w62_16 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1295_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1295_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1295_Out0_copy1296 :  std_logic_vector(2 downto 0);
signal bh793_w62_17 :  std_logic;
signal bh793_w63_15 :  std_logic;
signal bh793_w64_14 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1297_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1297_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1297_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1297_Out0_copy1298 :  std_logic_vector(2 downto 0);
signal bh793_w63_16 :  std_logic;
signal bh793_w64_15 :  std_logic;
signal bh793_w65_15 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1299_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1299_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1299_Out0_copy1300 :  std_logic_vector(1 downto 0);
signal bh793_w64_16 :  std_logic;
signal bh793_w65_16 :  std_logic;
signal Compressor_6_3_F200_uid1088_bh793_uid1301_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1301_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F200_uid1088_bh793_uid1301_Out0_copy1302 :  std_logic_vector(2 downto 0);
signal bh793_w65_17 :  std_logic;
signal bh793_w66_14 :  std_logic;
signal bh793_w67_13 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1303_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1303_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1303_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1303_Out0_copy1304 :  std_logic_vector(2 downto 0);
signal bh793_w66_15 :  std_logic;
signal bh793_w67_14 :  std_logic;
signal bh793_w68_14 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1305_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1305_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1305_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1305_Out0_copy1306 :  std_logic_vector(2 downto 0);
signal bh793_w67_15 :  std_logic;
signal bh793_w68_15 :  std_logic;
signal bh793_w69_12 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1307_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1307_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1307_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1307_Out0_copy1308 :  std_logic_vector(2 downto 0);
signal bh793_w68_16 :  std_logic;
signal bh793_w69_13 :  std_logic;
signal bh793_w70_13 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1309_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1309_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1309_Out0_copy1310 :  std_logic_vector(1 downto 0);
signal bh793_w69_14 :  std_logic;
signal bh793_w70_14 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1311_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1311_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1311_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1311_Out0_copy1312 :  std_logic_vector(2 downto 0);
signal bh793_w70_15 :  std_logic;
signal bh793_w71_14 :  std_logic;
signal bh793_w72_12 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1313_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1313_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1313_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1313_Out0_copy1314 :  std_logic_vector(2 downto 0);
signal bh793_w71_15 :  std_logic;
signal bh793_w72_13 :  std_logic;
signal bh793_w73_13 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1315_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1315_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1315_Out0_copy1316 :  std_logic_vector(1 downto 0);
signal bh793_w72_14 :  std_logic;
signal bh793_w73_14 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1317_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1317_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1317_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1317_Out0_copy1318 :  std_logic_vector(2 downto 0);
signal bh793_w73_15 :  std_logic;
signal bh793_w74_14 :  std_logic;
signal bh793_w75_12 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1319_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1319_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1319_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1319_Out0_copy1320 :  std_logic_vector(2 downto 0);
signal bh793_w74_15 :  std_logic;
signal bh793_w75_13 :  std_logic;
signal bh793_w76_13 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1321_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1321_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1321_Out0_copy1322 :  std_logic_vector(1 downto 0);
signal bh793_w75_14 :  std_logic;
signal bh793_w76_14 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1323_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1323_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1323_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1323_Out0_copy1324 :  std_logic_vector(2 downto 0);
signal bh793_w76_15 :  std_logic;
signal bh793_w77_12 :  std_logic;
signal bh793_w78_11 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1325_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1325_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1325_Out0_copy1326 :  std_logic_vector(1 downto 0);
signal bh793_w77_13 :  std_logic;
signal bh793_w78_12 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1327_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1327_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1327_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1327_Out0_copy1328 :  std_logic_vector(2 downto 0);
signal bh793_w78_13 :  std_logic;
signal bh793_w79_10 :  std_logic;
signal bh793_w80_12 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1329_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1329_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1329_Out0_copy1330 :  std_logic_vector(1 downto 0);
signal bh793_w79_11 :  std_logic;
signal bh793_w80_13 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1331_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1331_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1331_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1331_Out0_copy1332 :  std_logic_vector(2 downto 0);
signal bh793_w80_14 :  std_logic;
signal bh793_w81_11 :  std_logic;
signal bh793_w82_11 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1333_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1333_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1333_Out0_copy1334 :  std_logic_vector(1 downto 0);
signal bh793_w81_12 :  std_logic;
signal bh793_w82_12 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1335_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1335_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1335_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1335_Out0_copy1336 :  std_logic_vector(2 downto 0);
signal bh793_w82_13 :  std_logic;
signal bh793_w83_10 :  std_logic;
signal bh793_w84_9 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1337_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1337_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1337_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1337_Out0_copy1338 :  std_logic_vector(2 downto 0);
signal bh793_w83_11 :  std_logic;
signal bh793_w84_10 :  std_logic;
signal bh793_w85_10 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1339_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1339_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1339_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1339_Out0_copy1340 :  std_logic_vector(2 downto 0);
signal bh793_w85_11 :  std_logic;
signal bh793_w86_9 :  std_logic;
signal bh793_w87_9 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1341_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1341_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1341_Out0_copy1342 :  std_logic_vector(1 downto 0);
signal bh793_w86_10 :  std_logic;
signal bh793_w87_10 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1343_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1343_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1343_Out0_copy1344 :  std_logic_vector(1 downto 0);
signal bh793_w87_11 :  std_logic;
signal bh793_w88_10 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1345_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1345_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1345_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1345_Out0_copy1346 :  std_logic_vector(2 downto 0);
signal bh793_w88_11 :  std_logic;
signal bh793_w89_9 :  std_logic;
signal bh793_w90_9 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1347_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1347_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1347_Out0_copy1348 :  std_logic_vector(1 downto 0);
signal bh793_w89_10 :  std_logic;
signal bh793_w90_10 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1349_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1349_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1349_Out0_copy1350 :  std_logic_vector(1 downto 0);
signal bh793_w90_11 :  std_logic;
signal bh793_w91_10 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1351_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1351_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1351_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1351_Out0_copy1352 :  std_logic_vector(2 downto 0);
signal bh793_w91_11 :  std_logic;
signal bh793_w92_9 :  std_logic;
signal bh793_w93_9 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1353_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1353_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1353_Out0_copy1354 :  std_logic_vector(1 downto 0);
signal bh793_w92_10 :  std_logic;
signal bh793_w93_10 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1355_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1355_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1355_Out0_copy1356 :  std_logic_vector(1 downto 0);
signal bh793_w93_11 :  std_logic;
signal bh793_w94_10 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1357_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1357_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1357_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1357_Out0_copy1358 :  std_logic_vector(2 downto 0);
signal bh793_w94_11 :  std_logic;
signal bh793_w95_9 :  std_logic;
signal bh793_w96_9 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1359_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1359_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1359_Out0_copy1360 :  std_logic_vector(1 downto 0);
signal bh793_w95_10 :  std_logic;
signal bh793_w96_10 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1361_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1361_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1361_Out0_copy1362 :  std_logic_vector(1 downto 0);
signal bh793_w96_11 :  std_logic;
signal bh793_w97_10 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1363_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1363_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1363_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1363_Out0_copy1364 :  std_logic_vector(2 downto 0);
signal bh793_w97_11 :  std_logic;
signal bh793_w98_9 :  std_logic;
signal bh793_w99_9 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1365_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1365_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1365_Out0_copy1366 :  std_logic_vector(1 downto 0);
signal bh793_w98_10 :  std_logic;
signal bh793_w99_10 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1367_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1367_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1367_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1367_Out0_copy1368 :  std_logic_vector(2 downto 0);
signal bh793_w99_11 :  std_logic;
signal bh793_w100_9 :  std_logic;
signal bh793_w101_6 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1369_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1369_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1369_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1369_Out0_copy1370 :  std_logic_vector(2 downto 0);
signal bh793_w101_7 :  std_logic;
signal bh793_w102_7 :  std_logic;
signal bh793_w103_3 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1371_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1371_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1371_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1371_Out0_copy1372 :  std_logic_vector(2 downto 0);
signal bh793_w103_4 :  std_logic;
signal bh793_w104_2 :  std_logic;
signal bh793_w105_1 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1373_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1373_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1373_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1373_Out0_copy1374 :  std_logic_vector(2 downto 0);
signal bh793_w21_6 :  std_logic;
signal bh793_w22_4 :  std_logic;
signal bh793_w23_6 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1375_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1375_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1375_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1375_Out0_copy1376 :  std_logic_vector(2 downto 0);
signal bh793_w23_7 :  std_logic;
signal bh793_w24_6 :  std_logic;
signal bh793_w25_6 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1377_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1377_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1377_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1377_Out0_copy1378 :  std_logic_vector(2 downto 0);
signal bh793_w25_7 :  std_logic;
signal bh793_w26_6 :  std_logic;
signal bh793_w27_6 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1379_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1379_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1379_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1379_Out0_copy1380 :  std_logic_vector(2 downto 0);
signal bh793_w27_7 :  std_logic;
signal bh793_w28_6 :  std_logic;
signal bh793_w29_6 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1381_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1381_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1381_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1381_Out0_copy1382 :  std_logic_vector(2 downto 0);
signal bh793_w29_7 :  std_logic;
signal bh793_w30_6 :  std_logic;
signal bh793_w31_6 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1383_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1383_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1383_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1383_Out0_copy1384 :  std_logic_vector(2 downto 0);
signal bh793_w31_7 :  std_logic;
signal bh793_w32_6 :  std_logic;
signal bh793_w33_6 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1385_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1385_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1385_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1385_Out0_copy1386 :  std_logic_vector(2 downto 0);
signal bh793_w33_7 :  std_logic;
signal bh793_w34_7 :  std_logic;
signal bh793_w35_8 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1387_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1387_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1387_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1387_Out0_copy1388 :  std_logic_vector(2 downto 0);
signal bh793_w35_9 :  std_logic;
signal bh793_w36_9 :  std_logic;
signal bh793_w37_7 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1389_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1389_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1389_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1389_Out0_copy1390 :  std_logic_vector(2 downto 0);
signal bh793_w38_9 :  std_logic;
signal bh793_w39_7 :  std_logic;
signal bh793_w40_9 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1391_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1391_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1391_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1391_Out0_copy1392 :  std_logic_vector(2 downto 0);
signal bh793_w40_10 :  std_logic;
signal bh793_w41_7 :  std_logic;
signal bh793_w42_9 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1393_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1393_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1393_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1393_Out0_copy1394 :  std_logic_vector(2 downto 0);
signal bh793_w42_10 :  std_logic;
signal bh793_w43_7 :  std_logic;
signal bh793_w44_9 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1395_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1395_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1395_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1395_Out0_copy1396 :  std_logic_vector(2 downto 0);
signal bh793_w44_10 :  std_logic;
signal bh793_w45_7 :  std_logic;
signal bh793_w46_9 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1397_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1397_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1397_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1397_Out0_copy1398 :  std_logic_vector(2 downto 0);
signal bh793_w46_10 :  std_logic;
signal bh793_w47_7 :  std_logic;
signal bh793_w48_10 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1399_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1399_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1399_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1399_Out0_copy1400 :  std_logic_vector(2 downto 0);
signal bh793_w48_11 :  std_logic;
signal bh793_w49_9 :  std_logic;
signal bh793_w50_12 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1401_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1401_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1401_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1401_Out0_copy1402 :  std_logic_vector(2 downto 0);
signal bh793_w50_13 :  std_logic;
signal bh793_w51_12 :  std_logic;
signal bh793_w52_16 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1403_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1403_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1403_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1403_Out0_copy1404 :  std_logic_vector(2 downto 0);
signal bh793_w52_17 :  std_logic;
signal bh793_w53_15 :  std_logic;
signal bh793_w54_18 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1405_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1405_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1405_Out0_copy1406 :  std_logic_vector(1 downto 0);
signal bh793_w54_19 :  std_logic;
signal bh793_w55_17 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1407_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1407_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1407_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1407_Out0_copy1408 :  std_logic_vector(2 downto 0);
signal bh793_w55_18 :  std_logic;
signal bh793_w56_18 :  std_logic;
signal bh793_w57_17 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1409_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1409_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1409_Out0_copy1410 :  std_logic_vector(1 downto 0);
signal bh793_w56_19 :  std_logic;
signal bh793_w57_18 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1411_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1411_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1411_Out0_copy1412 :  std_logic_vector(1 downto 0);
signal bh793_w57_19 :  std_logic;
signal bh793_w58_17 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1413_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1413_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1413_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1413_Out0_copy1414 :  std_logic_vector(2 downto 0);
signal bh793_w58_18 :  std_logic;
signal bh793_w59_18 :  std_logic;
signal bh793_w60_17 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1415_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1415_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1415_Out0_copy1416 :  std_logic_vector(1 downto 0);
signal bh793_w59_19 :  std_logic;
signal bh793_w60_18 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1417_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1417_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1417_Out0_copy1418 :  std_logic_vector(1 downto 0);
signal bh793_w60_19 :  std_logic;
signal bh793_w61_17 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1419_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1419_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1419_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1419_Out0_copy1420 :  std_logic_vector(2 downto 0);
signal bh793_w61_18 :  std_logic;
signal bh793_w62_18 :  std_logic;
signal bh793_w63_17 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1421_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1421_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1421_Out0_copy1422 :  std_logic_vector(1 downto 0);
signal bh793_w62_19 :  std_logic;
signal bh793_w63_18 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1423_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1423_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1423_Out0_copy1424 :  std_logic_vector(1 downto 0);
signal bh793_w63_19 :  std_logic;
signal bh793_w64_17 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1425_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1425_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1425_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1425_Out0_copy1426 :  std_logic_vector(2 downto 0);
signal bh793_w64_18 :  std_logic;
signal bh793_w65_18 :  std_logic;
signal bh793_w66_16 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1427_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1427_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1427_Out0_copy1428 :  std_logic_vector(1 downto 0);
signal bh793_w65_19 :  std_logic;
signal bh793_w66_17 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1429_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1429_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1429_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1429_Out0_copy1430 :  std_logic_vector(2 downto 0);
signal bh793_w66_18 :  std_logic;
signal bh793_w67_16 :  std_logic;
signal bh793_w68_17 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1431_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1431_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1431_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1431_Out0_copy1432 :  std_logic_vector(2 downto 0);
signal bh793_w68_18 :  std_logic;
signal bh793_w69_15 :  std_logic;
signal bh793_w70_16 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1433_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1433_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1433_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1433_Out0_copy1434 :  std_logic_vector(2 downto 0);
signal bh793_w70_17 :  std_logic;
signal bh793_w71_16 :  std_logic;
signal bh793_w72_15 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1435_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1435_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1435_Out0_copy1436 :  std_logic_vector(1 downto 0);
signal bh793_w72_16 :  std_logic;
signal bh793_w73_16 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1437_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1437_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1437_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1437_Out0_copy1438 :  std_logic_vector(2 downto 0);
signal bh793_w73_17 :  std_logic;
signal bh793_w74_16 :  std_logic;
signal bh793_w75_15 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1439_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1439_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1439_Out0_copy1440 :  std_logic_vector(1 downto 0);
signal bh793_w75_16 :  std_logic;
signal bh793_w76_16 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1441_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1441_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1441_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1441_Out0_copy1442 :  std_logic_vector(2 downto 0);
signal bh793_w76_17 :  std_logic;
signal bh793_w77_14 :  std_logic;
signal bh793_w78_14 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1443_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1443_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1443_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1443_Out0_copy1444 :  std_logic_vector(2 downto 0);
signal bh793_w78_15 :  std_logic;
signal bh793_w79_12 :  std_logic;
signal bh793_w80_15 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1445_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1445_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1445_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1445_Out0_copy1446 :  std_logic_vector(2 downto 0);
signal bh793_w80_16 :  std_logic;
signal bh793_w81_13 :  std_logic;
signal bh793_w82_14 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1447_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1447_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1447_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1447_Out0_copy1448 :  std_logic_vector(2 downto 0);
signal bh793_w82_15 :  std_logic;
signal bh793_w83_12 :  std_logic;
signal bh793_w84_11 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1449_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1449_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1449_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1449_Out0_copy1450 :  std_logic_vector(2 downto 0);
signal bh793_w84_12 :  std_logic;
signal bh793_w85_12 :  std_logic;
signal bh793_w86_11 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1451_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1451_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1451_Out0_copy1452 :  std_logic_vector(1 downto 0);
signal bh793_w86_12 :  std_logic;
signal bh793_w87_12 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1453_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1453_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1453_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1453_Out0_copy1454 :  std_logic_vector(2 downto 0);
signal bh793_w87_13 :  std_logic;
signal bh793_w88_12 :  std_logic;
signal bh793_w89_11 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1455_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1455_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1455_Out0_copy1456 :  std_logic_vector(1 downto 0);
signal bh793_w89_12 :  std_logic;
signal bh793_w90_12 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1457_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1457_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1457_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1457_Out0_copy1458 :  std_logic_vector(2 downto 0);
signal bh793_w90_13 :  std_logic;
signal bh793_w91_12 :  std_logic;
signal bh793_w92_11 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1459_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1459_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1459_Out0_copy1460 :  std_logic_vector(1 downto 0);
signal bh793_w92_12 :  std_logic;
signal bh793_w93_12 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1461_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1461_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1461_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1461_Out0_copy1462 :  std_logic_vector(2 downto 0);
signal bh793_w93_13 :  std_logic;
signal bh793_w94_12 :  std_logic;
signal bh793_w95_11 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1463_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1463_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1463_Out0_copy1464 :  std_logic_vector(1 downto 0);
signal bh793_w95_12 :  std_logic;
signal bh793_w96_12 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1465_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1465_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1465_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1465_Out0_copy1466 :  std_logic_vector(2 downto 0);
signal bh793_w96_13 :  std_logic;
signal bh793_w97_12 :  std_logic;
signal bh793_w98_11 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1467_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1467_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1467_Out0_copy1468 :  std_logic_vector(1 downto 0);
signal bh793_w98_12 :  std_logic;
signal bh793_w99_12 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1469_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1469_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1469_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1469_Out0_copy1470 :  std_logic_vector(2 downto 0);
signal bh793_w99_13 :  std_logic;
signal bh793_w100_10 :  std_logic;
signal bh793_w101_8 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1471_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1471_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1471_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1471_Out0_copy1472 :  std_logic_vector(2 downto 0);
signal bh793_w101_9 :  std_logic;
signal bh793_w102_8 :  std_logic;
signal bh793_w103_5 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1473_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1473_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1473_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1473_Out0_copy1474 :  std_logic_vector(2 downto 0);
signal bh793_w103_6 :  std_logic;
signal bh793_w104_3 :  std_logic;
signal bh793_w105_2 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1475_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1475_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1475_Out0_copy1476 :  std_logic_vector(1 downto 0);
signal bh793_w105_3 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1477_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1477_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1477_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1477_Out0_copy1478 :  std_logic_vector(2 downto 0);
signal bh793_w23_8 :  std_logic;
signal bh793_w24_7 :  std_logic;
signal bh793_w25_8 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1479_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1479_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1479_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1479_Out0_copy1480 :  std_logic_vector(2 downto 0);
signal bh793_w25_9 :  std_logic;
signal bh793_w26_7 :  std_logic;
signal bh793_w27_8 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1481_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1481_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1481_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1481_Out0_copy1482 :  std_logic_vector(2 downto 0);
signal bh793_w27_9 :  std_logic;
signal bh793_w28_7 :  std_logic;
signal bh793_w29_8 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1483_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1483_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1483_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1483_Out0_copy1484 :  std_logic_vector(2 downto 0);
signal bh793_w29_9 :  std_logic;
signal bh793_w30_7 :  std_logic;
signal bh793_w31_8 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1485_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1485_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1485_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1485_Out0_copy1486 :  std_logic_vector(2 downto 0);
signal bh793_w31_9 :  std_logic;
signal bh793_w32_7 :  std_logic;
signal bh793_w33_8 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1487_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1487_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1487_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1487_Out0_copy1488 :  std_logic_vector(2 downto 0);
signal bh793_w33_9 :  std_logic;
signal bh793_w34_8 :  std_logic;
signal bh793_w35_10 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1489_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1489_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1489_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1489_Out0_copy1490 :  std_logic_vector(2 downto 0);
signal bh793_w35_11 :  std_logic;
signal bh793_w36_10 :  std_logic;
signal bh793_w37_8 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1491_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1491_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1491_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1491_Out0_copy1492 :  std_logic_vector(2 downto 0);
signal bh793_w37_9 :  std_logic;
signal bh793_w38_10 :  std_logic;
signal bh793_w39_8 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1493_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1493_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1493_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1493_Out0_copy1494 :  std_logic_vector(2 downto 0);
signal bh793_w40_11 :  std_logic;
signal bh793_w41_8 :  std_logic;
signal bh793_w42_11 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1495_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1495_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1495_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1495_Out0_copy1496 :  std_logic_vector(2 downto 0);
signal bh793_w42_12 :  std_logic;
signal bh793_w43_8 :  std_logic;
signal bh793_w44_11 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1497_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1497_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1497_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1497_Out0_copy1498 :  std_logic_vector(2 downto 0);
signal bh793_w44_12 :  std_logic;
signal bh793_w45_8 :  std_logic;
signal bh793_w46_11 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1499_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1499_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1499_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1499_Out0_copy1500 :  std_logic_vector(2 downto 0);
signal bh793_w46_12 :  std_logic;
signal bh793_w47_8 :  std_logic;
signal bh793_w48_12 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1501_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1501_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1501_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1501_Out0_copy1502 :  std_logic_vector(2 downto 0);
signal bh793_w48_13 :  std_logic;
signal bh793_w49_10 :  std_logic;
signal bh793_w50_14 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1503_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1503_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1503_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1503_Out0_copy1504 :  std_logic_vector(2 downto 0);
signal bh793_w50_15 :  std_logic;
signal bh793_w51_13 :  std_logic;
signal bh793_w52_18 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1505_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1505_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1505_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1505_Out0_copy1506 :  std_logic_vector(2 downto 0);
signal bh793_w52_19 :  std_logic;
signal bh793_w53_16 :  std_logic;
signal bh793_w54_20 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1507_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1507_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1507_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1507_Out0_copy1508 :  std_logic_vector(2 downto 0);
signal bh793_w54_21 :  std_logic;
signal bh793_w55_19 :  std_logic;
signal bh793_w56_20 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1509_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1509_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1509_Out0_copy1510 :  std_logic_vector(1 downto 0);
signal bh793_w56_21 :  std_logic;
signal bh793_w57_20 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1511_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1511_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1511_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1511_Out0_copy1512 :  std_logic_vector(2 downto 0);
signal bh793_w57_21 :  std_logic;
signal bh793_w58_19 :  std_logic;
signal bh793_w59_20 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1513_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1513_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1513_Out0_copy1514 :  std_logic_vector(1 downto 0);
signal bh793_w59_21 :  std_logic;
signal bh793_w60_20 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1515_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1515_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1515_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1515_Out0_copy1516 :  std_logic_vector(2 downto 0);
signal bh793_w60_21 :  std_logic;
signal bh793_w61_19 :  std_logic;
signal bh793_w62_20 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1517_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1517_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1517_Out0_copy1518 :  std_logic_vector(1 downto 0);
signal bh793_w62_21 :  std_logic;
signal bh793_w63_20 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1519_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1519_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1519_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1519_Out0_copy1520 :  std_logic_vector(2 downto 0);
signal bh793_w63_21 :  std_logic;
signal bh793_w64_19 :  std_logic;
signal bh793_w65_20 :  std_logic;
signal Compressor_3_2_F200_uid1040_bh793_uid1521_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1521_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F200_uid1040_bh793_uid1521_Out0_copy1522 :  std_logic_vector(1 downto 0);
signal bh793_w65_21 :  std_logic;
signal bh793_w66_19 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1523_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1523_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1523_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1523_Out0_copy1524 :  std_logic_vector(2 downto 0);
signal bh793_w66_20 :  std_logic;
signal bh793_w67_17 :  std_logic;
signal bh793_w68_19 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1525_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1525_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1525_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1525_Out0_copy1526 :  std_logic_vector(2 downto 0);
signal bh793_w68_20 :  std_logic;
signal bh793_w69_16 :  std_logic;
signal bh793_w70_18 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1527_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1527_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1527_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1527_Out0_copy1528 :  std_logic_vector(2 downto 0);
signal bh793_w70_19 :  std_logic;
signal bh793_w71_17 :  std_logic;
signal bh793_w72_17 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1529_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1529_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1529_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1529_Out0_copy1530 :  std_logic_vector(2 downto 0);
signal bh793_w72_18 :  std_logic;
signal bh793_w73_18 :  std_logic;
signal bh793_w74_17 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1531_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1531_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1531_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1531_Out0_copy1532 :  std_logic_vector(2 downto 0);
signal bh793_w74_18 :  std_logic;
signal bh793_w75_17 :  std_logic;
signal bh793_w76_18 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1533_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1533_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1533_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1533_Out0_copy1534 :  std_logic_vector(2 downto 0);
signal bh793_w76_19 :  std_logic;
signal bh793_w77_15 :  std_logic;
signal bh793_w78_16 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1535_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1535_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1535_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1535_Out0_copy1536 :  std_logic_vector(2 downto 0);
signal bh793_w78_17 :  std_logic;
signal bh793_w79_13 :  std_logic;
signal bh793_w80_17 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1537_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1537_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1537_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1537_Out0_copy1538 :  std_logic_vector(2 downto 0);
signal bh793_w80_18 :  std_logic;
signal bh793_w81_14 :  std_logic;
signal bh793_w82_16 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1539_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1539_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1539_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1539_Out0_copy1540 :  std_logic_vector(2 downto 0);
signal bh793_w82_17 :  std_logic;
signal bh793_w83_13 :  std_logic;
signal bh793_w84_13 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1541_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1541_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1541_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1541_Out0_copy1542 :  std_logic_vector(2 downto 0);
signal bh793_w84_14 :  std_logic;
signal bh793_w85_13 :  std_logic;
signal bh793_w86_13 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1543_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1543_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1543_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1543_Out0_copy1544 :  std_logic_vector(2 downto 0);
signal bh793_w86_14 :  std_logic;
signal bh793_w87_14 :  std_logic;
signal bh793_w88_13 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1545_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1545_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1545_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1545_Out0_copy1546 :  std_logic_vector(2 downto 0);
signal bh793_w89_13 :  std_logic;
signal bh793_w90_14 :  std_logic;
signal bh793_w91_13 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1547_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1547_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1547_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1547_Out0_copy1548 :  std_logic_vector(2 downto 0);
signal bh793_w92_13 :  std_logic;
signal bh793_w93_14 :  std_logic;
signal bh793_w94_13 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1549_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1549_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1549_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1549_Out0_copy1550 :  std_logic_vector(2 downto 0);
signal bh793_w95_13 :  std_logic;
signal bh793_w96_14 :  std_logic;
signal bh793_w97_13 :  std_logic;
signal Compressor_23_3_F200_uid1032_bh793_uid1551_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1551_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1551_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F200_uid1032_bh793_uid1551_Out0_copy1552 :  std_logic_vector(2 downto 0);
signal bh793_w98_13 :  std_logic;
signal bh793_w99_14 :  std_logic;
signal bh793_w100_11 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1553_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1553_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1553_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1553_Out0_copy1554 :  std_logic_vector(2 downto 0);
signal bh793_w101_10 :  std_logic;
signal bh793_w102_9 :  std_logic;
signal bh793_w103_7 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1555_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1555_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1555_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1555_Out0_copy1556 :  std_logic_vector(2 downto 0);
signal bh793_w103_8 :  std_logic;
signal bh793_w104_4 :  std_logic;
signal bh793_w105_4 :  std_logic;
signal Compressor_14_3_F200_uid1054_bh793_uid1557_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1557_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1557_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F200_uid1054_bh793_uid1557_Out0_copy1558 :  std_logic_vector(2 downto 0);
signal bh793_w105_5 :  std_logic;
signal tmp_bitheapResult_bh793_24 :  std_logic_vector(24 downto 0);
signal bitheapFinalAdd_bh793_In0 :  std_logic_vector(81 downto 0);
signal bitheapFinalAdd_bh793_In1 :  std_logic_vector(81 downto 0);
signal bitheapFinalAdd_bh793_Cin :  std_logic;
signal bitheapFinalAdd_bh793_Out :  std_logic_vector(81 downto 0);
signal bitheapResult_bh793 :  std_logic_vector(105 downto 0);
begin
   XX_m792 <= X ;
   YY_m792 <= Y ;
   tile_0_X <= X(16 downto 0);
   tile_0_Y <= Y(23 downto 0);
   tile_0_mult: DSPBlock_17x24_F200_uid795
      port map ( clk  => clk,
                 X => tile_0_X,
                 Y => tile_0_Y,
                 R => tile_0_output);

tile_0_filtered_output <= tile_0_output(40 downto 0);
   bh793_w0_0 <= tile_0_filtered_output(0);
   bh793_w1_0 <= tile_0_filtered_output(1);
   bh793_w2_0 <= tile_0_filtered_output(2);
   bh793_w3_0 <= tile_0_filtered_output(3);
   bh793_w4_0 <= tile_0_filtered_output(4);
   bh793_w5_0 <= tile_0_filtered_output(5);
   bh793_w6_0 <= tile_0_filtered_output(6);
   bh793_w7_0 <= tile_0_filtered_output(7);
   bh793_w8_0 <= tile_0_filtered_output(8);
   bh793_w9_0 <= tile_0_filtered_output(9);
   bh793_w10_0 <= tile_0_filtered_output(10);
   bh793_w11_0 <= tile_0_filtered_output(11);
   bh793_w12_0 <= tile_0_filtered_output(12);
   bh793_w13_0 <= tile_0_filtered_output(13);
   bh793_w14_0 <= tile_0_filtered_output(14);
   bh793_w15_0 <= tile_0_filtered_output(15);
   bh793_w16_0 <= tile_0_filtered_output(16);
   bh793_w17_0 <= tile_0_filtered_output(17);
   bh793_w18_0 <= tile_0_filtered_output(18);
   bh793_w19_0 <= tile_0_filtered_output(19);
   bh793_w20_0 <= tile_0_filtered_output(20);
   bh793_w21_0 <= tile_0_filtered_output(21);
   bh793_w22_0 <= tile_0_filtered_output(22);
   bh793_w23_0 <= tile_0_filtered_output(23);
   bh793_w24_0 <= tile_0_filtered_output(24);
   bh793_w25_0 <= tile_0_filtered_output(25);
   bh793_w26_0 <= tile_0_filtered_output(26);
   bh793_w27_0 <= tile_0_filtered_output(27);
   bh793_w28_0 <= tile_0_filtered_output(28);
   bh793_w29_0 <= tile_0_filtered_output(29);
   bh793_w30_0 <= tile_0_filtered_output(30);
   bh793_w31_0 <= tile_0_filtered_output(31);
   bh793_w32_0 <= tile_0_filtered_output(32);
   bh793_w33_0 <= tile_0_filtered_output(33);
   bh793_w34_0 <= tile_0_filtered_output(34);
   bh793_w35_0 <= tile_0_filtered_output(35);
   bh793_w36_0 <= tile_0_filtered_output(36);
   bh793_w37_0 <= tile_0_filtered_output(37);
   bh793_w38_0 <= tile_0_filtered_output(38);
   bh793_w39_0 <= tile_0_filtered_output(39);
   bh793_w40_0 <= tile_0_filtered_output(40);
   tile_1_X <= X(33 downto 17);
   tile_1_Y <= Y(23 downto 0);
   tile_1_mult: DSPBlock_17x24_F200_uid797
      port map ( clk  => clk,
                 X => tile_1_X,
                 Y => tile_1_Y,
                 R => tile_1_output);

tile_1_filtered_output <= tile_1_output(40 downto 0);
   bh793_w17_1 <= tile_1_filtered_output(0);
   bh793_w18_1 <= tile_1_filtered_output(1);
   bh793_w19_1 <= tile_1_filtered_output(2);
   bh793_w20_1 <= tile_1_filtered_output(3);
   bh793_w21_1 <= tile_1_filtered_output(4);
   bh793_w22_1 <= tile_1_filtered_output(5);
   bh793_w23_1 <= tile_1_filtered_output(6);
   bh793_w24_1 <= tile_1_filtered_output(7);
   bh793_w25_1 <= tile_1_filtered_output(8);
   bh793_w26_1 <= tile_1_filtered_output(9);
   bh793_w27_1 <= tile_1_filtered_output(10);
   bh793_w28_1 <= tile_1_filtered_output(11);
   bh793_w29_1 <= tile_1_filtered_output(12);
   bh793_w30_1 <= tile_1_filtered_output(13);
   bh793_w31_1 <= tile_1_filtered_output(14);
   bh793_w32_1 <= tile_1_filtered_output(15);
   bh793_w33_1 <= tile_1_filtered_output(16);
   bh793_w34_1 <= tile_1_filtered_output(17);
   bh793_w35_1 <= tile_1_filtered_output(18);
   bh793_w36_1 <= tile_1_filtered_output(19);
   bh793_w37_1 <= tile_1_filtered_output(20);
   bh793_w38_1 <= tile_1_filtered_output(21);
   bh793_w39_1 <= tile_1_filtered_output(22);
   bh793_w40_1 <= tile_1_filtered_output(23);
   bh793_w41_0 <= tile_1_filtered_output(24);
   bh793_w42_0 <= tile_1_filtered_output(25);
   bh793_w43_0 <= tile_1_filtered_output(26);
   bh793_w44_0 <= tile_1_filtered_output(27);
   bh793_w45_0 <= tile_1_filtered_output(28);
   bh793_w46_0 <= tile_1_filtered_output(29);
   bh793_w47_0 <= tile_1_filtered_output(30);
   bh793_w48_0 <= tile_1_filtered_output(31);
   bh793_w49_0 <= tile_1_filtered_output(32);
   bh793_w50_0 <= tile_1_filtered_output(33);
   bh793_w51_0 <= tile_1_filtered_output(34);
   bh793_w52_0 <= tile_1_filtered_output(35);
   bh793_w53_0 <= tile_1_filtered_output(36);
   bh793_w54_0 <= tile_1_filtered_output(37);
   bh793_w55_0 <= tile_1_filtered_output(38);
   bh793_w56_0 <= tile_1_filtered_output(39);
   bh793_w57_0 <= tile_1_filtered_output(40);
   tile_2_X <= X(50 downto 34);
   tile_2_Y <= Y(23 downto 0);
   tile_2_mult: DSPBlock_17x24_F200_uid799
      port map ( clk  => clk,
                 X => tile_2_X,
                 Y => tile_2_Y,
                 R => tile_2_output);

tile_2_filtered_output <= tile_2_output(40 downto 0);
   bh793_w34_2 <= tile_2_filtered_output(0);
   bh793_w35_2 <= tile_2_filtered_output(1);
   bh793_w36_2 <= tile_2_filtered_output(2);
   bh793_w37_2 <= tile_2_filtered_output(3);
   bh793_w38_2 <= tile_2_filtered_output(4);
   bh793_w39_2 <= tile_2_filtered_output(5);
   bh793_w40_2 <= tile_2_filtered_output(6);
   bh793_w41_1 <= tile_2_filtered_output(7);
   bh793_w42_1 <= tile_2_filtered_output(8);
   bh793_w43_1 <= tile_2_filtered_output(9);
   bh793_w44_1 <= tile_2_filtered_output(10);
   bh793_w45_1 <= tile_2_filtered_output(11);
   bh793_w46_1 <= tile_2_filtered_output(12);
   bh793_w47_1 <= tile_2_filtered_output(13);
   bh793_w48_1 <= tile_2_filtered_output(14);
   bh793_w49_1 <= tile_2_filtered_output(15);
   bh793_w50_1 <= tile_2_filtered_output(16);
   bh793_w51_1 <= tile_2_filtered_output(17);
   bh793_w52_1 <= tile_2_filtered_output(18);
   bh793_w53_1 <= tile_2_filtered_output(19);
   bh793_w54_1 <= tile_2_filtered_output(20);
   bh793_w55_1 <= tile_2_filtered_output(21);
   bh793_w56_1 <= tile_2_filtered_output(22);
   bh793_w57_1 <= tile_2_filtered_output(23);
   bh793_w58_0 <= tile_2_filtered_output(24);
   bh793_w59_0 <= tile_2_filtered_output(25);
   bh793_w60_0 <= tile_2_filtered_output(26);
   bh793_w61_0 <= tile_2_filtered_output(27);
   bh793_w62_0 <= tile_2_filtered_output(28);
   bh793_w63_0 <= tile_2_filtered_output(29);
   bh793_w64_0 <= tile_2_filtered_output(30);
   bh793_w65_0 <= tile_2_filtered_output(31);
   bh793_w66_0 <= tile_2_filtered_output(32);
   bh793_w67_0 <= tile_2_filtered_output(33);
   bh793_w68_0 <= tile_2_filtered_output(34);
   bh793_w69_0 <= tile_2_filtered_output(35);
   bh793_w70_0 <= tile_2_filtered_output(36);
   bh793_w71_0 <= tile_2_filtered_output(37);
   bh793_w72_0 <= tile_2_filtered_output(38);
   bh793_w73_0 <= tile_2_filtered_output(39);
   bh793_w74_0 <= tile_2_filtered_output(40);
   tile_3_X <= X(52 downto 51);
   tile_3_Y <= Y(23 downto 0);
   tile_3_mult: DSPBlock_2x24_F200_uid801
      port map ( clk  => clk,
                 X => tile_3_X,
                 Y => tile_3_Y,
                 R => tile_3_output);

tile_3_filtered_output <= tile_3_output(25 downto 0);
   bh793_w51_2 <= tile_3_filtered_output(0);
   bh793_w52_2 <= tile_3_filtered_output(1);
   bh793_w53_2 <= tile_3_filtered_output(2);
   bh793_w54_2 <= tile_3_filtered_output(3);
   bh793_w55_2 <= tile_3_filtered_output(4);
   bh793_w56_2 <= tile_3_filtered_output(5);
   bh793_w57_2 <= tile_3_filtered_output(6);
   bh793_w58_1 <= tile_3_filtered_output(7);
   bh793_w59_1 <= tile_3_filtered_output(8);
   bh793_w60_1 <= tile_3_filtered_output(9);
   bh793_w61_1 <= tile_3_filtered_output(10);
   bh793_w62_1 <= tile_3_filtered_output(11);
   bh793_w63_1 <= tile_3_filtered_output(12);
   bh793_w64_1 <= tile_3_filtered_output(13);
   bh793_w65_1 <= tile_3_filtered_output(14);
   bh793_w66_1 <= tile_3_filtered_output(15);
   bh793_w67_1 <= tile_3_filtered_output(16);
   bh793_w68_1 <= tile_3_filtered_output(17);
   bh793_w69_1 <= tile_3_filtered_output(18);
   bh793_w70_1 <= tile_3_filtered_output(19);
   bh793_w71_1 <= tile_3_filtered_output(20);
   bh793_w72_1 <= tile_3_filtered_output(21);
   bh793_w73_1 <= tile_3_filtered_output(22);
   bh793_w74_1 <= tile_3_filtered_output(23);
   bh793_w75_0 <= tile_3_filtered_output(24);
   bh793_w76_0 <= tile_3_filtered_output(25);
   tile_4_X <= X(16 downto 0);
   tile_4_Y <= Y(47 downto 24);
   tile_4_mult: DSPBlock_17x24_F200_uid803
      port map ( clk  => clk,
                 X => tile_4_X,
                 Y => tile_4_Y,
                 R => tile_4_output);

tile_4_filtered_output <= tile_4_output(40 downto 0);
   bh793_w24_2 <= tile_4_filtered_output(0);
   bh793_w25_2 <= tile_4_filtered_output(1);
   bh793_w26_2 <= tile_4_filtered_output(2);
   bh793_w27_2 <= tile_4_filtered_output(3);
   bh793_w28_2 <= tile_4_filtered_output(4);
   bh793_w29_2 <= tile_4_filtered_output(5);
   bh793_w30_2 <= tile_4_filtered_output(6);
   bh793_w31_2 <= tile_4_filtered_output(7);
   bh793_w32_2 <= tile_4_filtered_output(8);
   bh793_w33_2 <= tile_4_filtered_output(9);
   bh793_w34_3 <= tile_4_filtered_output(10);
   bh793_w35_3 <= tile_4_filtered_output(11);
   bh793_w36_3 <= tile_4_filtered_output(12);
   bh793_w37_3 <= tile_4_filtered_output(13);
   bh793_w38_3 <= tile_4_filtered_output(14);
   bh793_w39_3 <= tile_4_filtered_output(15);
   bh793_w40_3 <= tile_4_filtered_output(16);
   bh793_w41_2 <= tile_4_filtered_output(17);
   bh793_w42_2 <= tile_4_filtered_output(18);
   bh793_w43_2 <= tile_4_filtered_output(19);
   bh793_w44_2 <= tile_4_filtered_output(20);
   bh793_w45_2 <= tile_4_filtered_output(21);
   bh793_w46_2 <= tile_4_filtered_output(22);
   bh793_w47_2 <= tile_4_filtered_output(23);
   bh793_w48_2 <= tile_4_filtered_output(24);
   bh793_w49_2 <= tile_4_filtered_output(25);
   bh793_w50_2 <= tile_4_filtered_output(26);
   bh793_w51_3 <= tile_4_filtered_output(27);
   bh793_w52_3 <= tile_4_filtered_output(28);
   bh793_w53_3 <= tile_4_filtered_output(29);
   bh793_w54_3 <= tile_4_filtered_output(30);
   bh793_w55_3 <= tile_4_filtered_output(31);
   bh793_w56_3 <= tile_4_filtered_output(32);
   bh793_w57_3 <= tile_4_filtered_output(33);
   bh793_w58_2 <= tile_4_filtered_output(34);
   bh793_w59_2 <= tile_4_filtered_output(35);
   bh793_w60_2 <= tile_4_filtered_output(36);
   bh793_w61_2 <= tile_4_filtered_output(37);
   bh793_w62_2 <= tile_4_filtered_output(38);
   bh793_w63_2 <= tile_4_filtered_output(39);
   bh793_w64_2 <= tile_4_filtered_output(40);
   tile_5_X <= X(33 downto 17);
   tile_5_Y <= Y(47 downto 24);
   tile_5_mult: DSPBlock_17x24_F200_uid805
      port map ( clk  => clk,
                 X => tile_5_X,
                 Y => tile_5_Y,
                 R => tile_5_output);

tile_5_filtered_output <= tile_5_output(40 downto 0);
   bh793_w41_3 <= tile_5_filtered_output(0);
   bh793_w42_3 <= tile_5_filtered_output(1);
   bh793_w43_3 <= tile_5_filtered_output(2);
   bh793_w44_3 <= tile_5_filtered_output(3);
   bh793_w45_3 <= tile_5_filtered_output(4);
   bh793_w46_3 <= tile_5_filtered_output(5);
   bh793_w47_3 <= tile_5_filtered_output(6);
   bh793_w48_3 <= tile_5_filtered_output(7);
   bh793_w49_3 <= tile_5_filtered_output(8);
   bh793_w50_3 <= tile_5_filtered_output(9);
   bh793_w51_4 <= tile_5_filtered_output(10);
   bh793_w52_4 <= tile_5_filtered_output(11);
   bh793_w53_4 <= tile_5_filtered_output(12);
   bh793_w54_4 <= tile_5_filtered_output(13);
   bh793_w55_4 <= tile_5_filtered_output(14);
   bh793_w56_4 <= tile_5_filtered_output(15);
   bh793_w57_4 <= tile_5_filtered_output(16);
   bh793_w58_3 <= tile_5_filtered_output(17);
   bh793_w59_3 <= tile_5_filtered_output(18);
   bh793_w60_3 <= tile_5_filtered_output(19);
   bh793_w61_3 <= tile_5_filtered_output(20);
   bh793_w62_3 <= tile_5_filtered_output(21);
   bh793_w63_3 <= tile_5_filtered_output(22);
   bh793_w64_3 <= tile_5_filtered_output(23);
   bh793_w65_2 <= tile_5_filtered_output(24);
   bh793_w66_2 <= tile_5_filtered_output(25);
   bh793_w67_2 <= tile_5_filtered_output(26);
   bh793_w68_2 <= tile_5_filtered_output(27);
   bh793_w69_2 <= tile_5_filtered_output(28);
   bh793_w70_2 <= tile_5_filtered_output(29);
   bh793_w71_2 <= tile_5_filtered_output(30);
   bh793_w72_2 <= tile_5_filtered_output(31);
   bh793_w73_2 <= tile_5_filtered_output(32);
   bh793_w74_2 <= tile_5_filtered_output(33);
   bh793_w75_1 <= tile_5_filtered_output(34);
   bh793_w76_1 <= tile_5_filtered_output(35);
   bh793_w77_0 <= tile_5_filtered_output(36);
   bh793_w78_0 <= tile_5_filtered_output(37);
   bh793_w79_0 <= tile_5_filtered_output(38);
   bh793_w80_0 <= tile_5_filtered_output(39);
   bh793_w81_0 <= tile_5_filtered_output(40);
   tile_6_X <= X(50 downto 34);
   tile_6_Y <= Y(47 downto 24);
   tile_6_mult: DSPBlock_17x24_F200_uid807
      port map ( clk  => clk,
                 X => tile_6_X,
                 Y => tile_6_Y,
                 R => tile_6_output);

tile_6_filtered_output <= tile_6_output(40 downto 0);
   bh793_w58_4 <= tile_6_filtered_output(0);
   bh793_w59_4 <= tile_6_filtered_output(1);
   bh793_w60_4 <= tile_6_filtered_output(2);
   bh793_w61_4 <= tile_6_filtered_output(3);
   bh793_w62_4 <= tile_6_filtered_output(4);
   bh793_w63_4 <= tile_6_filtered_output(5);
   bh793_w64_4 <= tile_6_filtered_output(6);
   bh793_w65_3 <= tile_6_filtered_output(7);
   bh793_w66_3 <= tile_6_filtered_output(8);
   bh793_w67_3 <= tile_6_filtered_output(9);
   bh793_w68_3 <= tile_6_filtered_output(10);
   bh793_w69_3 <= tile_6_filtered_output(11);
   bh793_w70_3 <= tile_6_filtered_output(12);
   bh793_w71_3 <= tile_6_filtered_output(13);
   bh793_w72_3 <= tile_6_filtered_output(14);
   bh793_w73_3 <= tile_6_filtered_output(15);
   bh793_w74_3 <= tile_6_filtered_output(16);
   bh793_w75_2 <= tile_6_filtered_output(17);
   bh793_w76_2 <= tile_6_filtered_output(18);
   bh793_w77_1 <= tile_6_filtered_output(19);
   bh793_w78_1 <= tile_6_filtered_output(20);
   bh793_w79_1 <= tile_6_filtered_output(21);
   bh793_w80_1 <= tile_6_filtered_output(22);
   bh793_w81_1 <= tile_6_filtered_output(23);
   bh793_w82_0 <= tile_6_filtered_output(24);
   bh793_w83_0 <= tile_6_filtered_output(25);
   bh793_w84_0 <= tile_6_filtered_output(26);
   bh793_w85_0 <= tile_6_filtered_output(27);
   bh793_w86_0 <= tile_6_filtered_output(28);
   bh793_w87_0 <= tile_6_filtered_output(29);
   bh793_w88_0 <= tile_6_filtered_output(30);
   bh793_w89_0 <= tile_6_filtered_output(31);
   bh793_w90_0 <= tile_6_filtered_output(32);
   bh793_w91_0 <= tile_6_filtered_output(33);
   bh793_w92_0 <= tile_6_filtered_output(34);
   bh793_w93_0 <= tile_6_filtered_output(35);
   bh793_w94_0 <= tile_6_filtered_output(36);
   bh793_w95_0 <= tile_6_filtered_output(37);
   bh793_w96_0 <= tile_6_filtered_output(38);
   bh793_w97_0 <= tile_6_filtered_output(39);
   bh793_w98_0 <= tile_6_filtered_output(40);
   tile_7_X <= X(52 downto 51);
   tile_7_Y <= Y(47 downto 24);
   tile_7_mult: DSPBlock_2x24_F200_uid809
      port map ( clk  => clk,
                 X => tile_7_X,
                 Y => tile_7_Y,
                 R => tile_7_output);

tile_7_filtered_output <= tile_7_output(25 downto 0);
   bh793_w75_3 <= tile_7_filtered_output(0);
   bh793_w76_3 <= tile_7_filtered_output(1);
   bh793_w77_2 <= tile_7_filtered_output(2);
   bh793_w78_2 <= tile_7_filtered_output(3);
   bh793_w79_2 <= tile_7_filtered_output(4);
   bh793_w80_2 <= tile_7_filtered_output(5);
   bh793_w81_2 <= tile_7_filtered_output(6);
   bh793_w82_1 <= tile_7_filtered_output(7);
   bh793_w83_1 <= tile_7_filtered_output(8);
   bh793_w84_1 <= tile_7_filtered_output(9);
   bh793_w85_1 <= tile_7_filtered_output(10);
   bh793_w86_1 <= tile_7_filtered_output(11);
   bh793_w87_1 <= tile_7_filtered_output(12);
   bh793_w88_1 <= tile_7_filtered_output(13);
   bh793_w89_1 <= tile_7_filtered_output(14);
   bh793_w90_1 <= tile_7_filtered_output(15);
   bh793_w91_1 <= tile_7_filtered_output(16);
   bh793_w92_1 <= tile_7_filtered_output(17);
   bh793_w93_1 <= tile_7_filtered_output(18);
   bh793_w94_1 <= tile_7_filtered_output(19);
   bh793_w95_1 <= tile_7_filtered_output(20);
   bh793_w96_1 <= tile_7_filtered_output(21);
   bh793_w97_1 <= tile_7_filtered_output(22);
   bh793_w98_1 <= tile_7_filtered_output(23);
   bh793_w99_0 <= tile_7_filtered_output(24);
   bh793_w100_0 <= tile_7_filtered_output(25);
   tile_8_X <= X(16 downto 16);
   tile_8_Y <= Y(52 downto 52);
   tile_8_mult: IntMultiplierLUT_1x1_F200_uid811
      port map ( clk  => clk,
                 X => tile_8_X,
                 Y => tile_8_Y,
                 R => tile_8_output);

tile_8_filtered_output <= tile_8_output(0 downto 0);
   bh793_w68_4 <= tile_8_filtered_output(0);
   tile_9_X <= X(15 downto 12);
   tile_9_Y <= Y(52 downto 52);
   tile_9_mult: IntMultiplierLUT_4x1_F200_uid813
      port map ( clk  => clk,
                 X => tile_9_X,
                 Y => tile_9_Y,
                 R => tile_9_output);

tile_9_filtered_output <= tile_9_output(3 downto 0);
   bh793_w64_5 <= tile_9_filtered_output(0);
   bh793_w65_4 <= tile_9_filtered_output(1);
   bh793_w66_4 <= tile_9_filtered_output(2);
   bh793_w67_4 <= tile_9_filtered_output(3);
   tile_10_X <= X(11 downto 8);
   tile_10_Y <= Y(52 downto 52);
   tile_10_mult: IntMultiplierLUT_4x1_F200_uid815
      port map ( clk  => clk,
                 X => tile_10_X,
                 Y => tile_10_Y,
                 R => tile_10_output);

tile_10_filtered_output <= tile_10_output(3 downto 0);
   bh793_w60_5 <= tile_10_filtered_output(0);
   bh793_w61_5 <= tile_10_filtered_output(1);
   bh793_w62_5 <= tile_10_filtered_output(2);
   bh793_w63_5 <= tile_10_filtered_output(3);
   tile_11_X <= X(7 downto 4);
   tile_11_Y <= Y(52 downto 52);
   tile_11_mult: IntMultiplierLUT_4x1_F200_uid817
      port map ( clk  => clk,
                 X => tile_11_X,
                 Y => tile_11_Y,
                 R => tile_11_output);

tile_11_filtered_output <= tile_11_output(3 downto 0);
   bh793_w56_5 <= tile_11_filtered_output(0);
   bh793_w57_5 <= tile_11_filtered_output(1);
   bh793_w58_5 <= tile_11_filtered_output(2);
   bh793_w59_5 <= tile_11_filtered_output(3);
   tile_12_X <= X(3 downto 0);
   tile_12_Y <= Y(52 downto 52);
   tile_12_mult: IntMultiplierLUT_4x1_F200_uid819
      port map ( clk  => clk,
                 X => tile_12_X,
                 Y => tile_12_Y,
                 R => tile_12_output);

tile_12_filtered_output <= tile_12_output(3 downto 0);
   bh793_w52_5 <= tile_12_filtered_output(0);
   bh793_w53_5 <= tile_12_filtered_output(1);
   bh793_w54_5 <= tile_12_filtered_output(2);
   bh793_w55_5 <= tile_12_filtered_output(3);
   tile_13_X <= X(16 downto 15);
   tile_13_Y <= Y(51 downto 50);
   tile_13_mult: IntMultiplierLUT_2x2_F200_uid821
      port map ( clk  => clk,
                 X => tile_13_X,
                 Y => tile_13_Y,
                 R => tile_13_output);

tile_13_filtered_output <= tile_13_output(3 downto 0);
   bh793_w65_5 <= tile_13_filtered_output(0);
   bh793_w66_5 <= tile_13_filtered_output(1);
   bh793_w67_5 <= tile_13_filtered_output(2);
   bh793_w68_5 <= tile_13_filtered_output(3);
   tile_14_X <= X(14 downto 12);
   tile_14_Y <= Y(51 downto 50);
   tile_14_mult: IntMultiplierLUT_3x2_F200_uid826
      port map ( clk  => clk,
                 X => tile_14_X,
                 Y => tile_14_Y,
                 R => tile_14_output);

tile_14_filtered_output <= tile_14_output(4 downto 0);
   bh793_w62_6 <= tile_14_filtered_output(0);
   bh793_w63_6 <= tile_14_filtered_output(1);
   bh793_w64_6 <= tile_14_filtered_output(2);
   bh793_w65_6 <= tile_14_filtered_output(3);
   bh793_w66_6 <= tile_14_filtered_output(4);
   tile_15_X <= X(11 downto 9);
   tile_15_Y <= Y(51 downto 50);
   tile_15_mult: IntMultiplierLUT_3x2_F200_uid831
      port map ( clk  => clk,
                 X => tile_15_X,
                 Y => tile_15_Y,
                 R => tile_15_output);

tile_15_filtered_output <= tile_15_output(4 downto 0);
   bh793_w59_6 <= tile_15_filtered_output(0);
   bh793_w60_6 <= tile_15_filtered_output(1);
   bh793_w61_6 <= tile_15_filtered_output(2);
   bh793_w62_7 <= tile_15_filtered_output(3);
   bh793_w63_7 <= tile_15_filtered_output(4);
   tile_16_X <= X(8 downto 6);
   tile_16_Y <= Y(51 downto 50);
   tile_16_mult: IntMultiplierLUT_3x2_F200_uid836
      port map ( clk  => clk,
                 X => tile_16_X,
                 Y => tile_16_Y,
                 R => tile_16_output);

tile_16_filtered_output <= tile_16_output(4 downto 0);
   bh793_w56_6 <= tile_16_filtered_output(0);
   bh793_w57_6 <= tile_16_filtered_output(1);
   bh793_w58_6 <= tile_16_filtered_output(2);
   bh793_w59_7 <= tile_16_filtered_output(3);
   bh793_w60_7 <= tile_16_filtered_output(4);
   tile_17_X <= X(5 downto 3);
   tile_17_Y <= Y(51 downto 50);
   tile_17_mult: IntMultiplierLUT_3x2_F200_uid841
      port map ( clk  => clk,
                 X => tile_17_X,
                 Y => tile_17_Y,
                 R => tile_17_output);

tile_17_filtered_output <= tile_17_output(4 downto 0);
   bh793_w53_6 <= tile_17_filtered_output(0);
   bh793_w54_6 <= tile_17_filtered_output(1);
   bh793_w55_6 <= tile_17_filtered_output(2);
   bh793_w56_7 <= tile_17_filtered_output(3);
   bh793_w57_7 <= tile_17_filtered_output(4);
   tile_18_X <= X(2 downto 0);
   tile_18_Y <= Y(51 downto 50);
   tile_18_mult: IntMultiplierLUT_3x2_F200_uid846
      port map ( clk  => clk,
                 X => tile_18_X,
                 Y => tile_18_Y,
                 R => tile_18_output);

tile_18_filtered_output <= tile_18_output(4 downto 0);
   bh793_w50_4 <= tile_18_filtered_output(0);
   bh793_w51_5 <= tile_18_filtered_output(1);
   bh793_w52_6 <= tile_18_filtered_output(2);
   bh793_w53_7 <= tile_18_filtered_output(3);
   bh793_w54_7 <= tile_18_filtered_output(4);
   tile_19_X <= X(16 downto 15);
   tile_19_Y <= Y(49 downto 48);
   tile_19_mult: IntMultiplierLUT_2x2_F200_uid851
      port map ( clk  => clk,
                 X => tile_19_X,
                 Y => tile_19_Y,
                 R => tile_19_output);

tile_19_filtered_output <= tile_19_output(3 downto 0);
   bh793_w63_8 <= tile_19_filtered_output(0);
   bh793_w64_7 <= tile_19_filtered_output(1);
   bh793_w65_7 <= tile_19_filtered_output(2);
   bh793_w66_7 <= tile_19_filtered_output(3);
   tile_20_X <= X(14 downto 12);
   tile_20_Y <= Y(49 downto 48);
   tile_20_mult: IntMultiplierLUT_3x2_F200_uid856
      port map ( clk  => clk,
                 X => tile_20_X,
                 Y => tile_20_Y,
                 R => tile_20_output);

tile_20_filtered_output <= tile_20_output(4 downto 0);
   bh793_w60_8 <= tile_20_filtered_output(0);
   bh793_w61_7 <= tile_20_filtered_output(1);
   bh793_w62_8 <= tile_20_filtered_output(2);
   bh793_w63_9 <= tile_20_filtered_output(3);
   bh793_w64_8 <= tile_20_filtered_output(4);
   tile_21_X <= X(11 downto 9);
   tile_21_Y <= Y(49 downto 48);
   tile_21_mult: IntMultiplierLUT_3x2_F200_uid861
      port map ( clk  => clk,
                 X => tile_21_X,
                 Y => tile_21_Y,
                 R => tile_21_output);

tile_21_filtered_output <= tile_21_output(4 downto 0);
   bh793_w57_8 <= tile_21_filtered_output(0);
   bh793_w58_7 <= tile_21_filtered_output(1);
   bh793_w59_8 <= tile_21_filtered_output(2);
   bh793_w60_9 <= tile_21_filtered_output(3);
   bh793_w61_8 <= tile_21_filtered_output(4);
   tile_22_X <= X(8 downto 6);
   tile_22_Y <= Y(49 downto 48);
   tile_22_mult: IntMultiplierLUT_3x2_F200_uid866
      port map ( clk  => clk,
                 X => tile_22_X,
                 Y => tile_22_Y,
                 R => tile_22_output);

tile_22_filtered_output <= tile_22_output(4 downto 0);
   bh793_w54_8 <= tile_22_filtered_output(0);
   bh793_w55_7 <= tile_22_filtered_output(1);
   bh793_w56_8 <= tile_22_filtered_output(2);
   bh793_w57_9 <= tile_22_filtered_output(3);
   bh793_w58_8 <= tile_22_filtered_output(4);
   tile_23_X <= X(5 downto 3);
   tile_23_Y <= Y(49 downto 48);
   tile_23_mult: IntMultiplierLUT_3x2_F200_uid871
      port map ( clk  => clk,
                 X => tile_23_X,
                 Y => tile_23_Y,
                 R => tile_23_output);

tile_23_filtered_output <= tile_23_output(4 downto 0);
   bh793_w51_6 <= tile_23_filtered_output(0);
   bh793_w52_7 <= tile_23_filtered_output(1);
   bh793_w53_8 <= tile_23_filtered_output(2);
   bh793_w54_9 <= tile_23_filtered_output(3);
   bh793_w55_8 <= tile_23_filtered_output(4);
   tile_24_X <= X(2 downto 0);
   tile_24_Y <= Y(49 downto 48);
   tile_24_mult: IntMultiplierLUT_3x2_F200_uid876
      port map ( clk  => clk,
                 X => tile_24_X,
                 Y => tile_24_Y,
                 R => tile_24_output);

tile_24_filtered_output <= tile_24_output(4 downto 0);
   bh793_w48_4 <= tile_24_filtered_output(0);
   bh793_w49_4 <= tile_24_filtered_output(1);
   bh793_w50_5 <= tile_24_filtered_output(2);
   bh793_w51_7 <= tile_24_filtered_output(3);
   bh793_w52_8 <= tile_24_filtered_output(4);
   tile_25_X <= X(33 downto 33);
   tile_25_Y <= Y(52 downto 52);
   tile_25_mult: IntMultiplierLUT_1x1_F200_uid881
      port map ( clk  => clk,
                 X => tile_25_X,
                 Y => tile_25_Y,
                 R => tile_25_output);

tile_25_filtered_output <= tile_25_output(0 downto 0);
   bh793_w85_2 <= tile_25_filtered_output(0);
   tile_26_X <= X(32 downto 29);
   tile_26_Y <= Y(52 downto 52);
   tile_26_mult: IntMultiplierLUT_4x1_F200_uid883
      port map ( clk  => clk,
                 X => tile_26_X,
                 Y => tile_26_Y,
                 R => tile_26_output);

tile_26_filtered_output <= tile_26_output(3 downto 0);
   bh793_w81_3 <= tile_26_filtered_output(0);
   bh793_w82_2 <= tile_26_filtered_output(1);
   bh793_w83_2 <= tile_26_filtered_output(2);
   bh793_w84_2 <= tile_26_filtered_output(3);
   tile_27_X <= X(28 downto 25);
   tile_27_Y <= Y(52 downto 52);
   tile_27_mult: IntMultiplierLUT_4x1_F200_uid885
      port map ( clk  => clk,
                 X => tile_27_X,
                 Y => tile_27_Y,
                 R => tile_27_output);

tile_27_filtered_output <= tile_27_output(3 downto 0);
   bh793_w77_3 <= tile_27_filtered_output(0);
   bh793_w78_3 <= tile_27_filtered_output(1);
   bh793_w79_3 <= tile_27_filtered_output(2);
   bh793_w80_3 <= tile_27_filtered_output(3);
   tile_28_X <= X(24 downto 21);
   tile_28_Y <= Y(52 downto 52);
   tile_28_mult: IntMultiplierLUT_4x1_F200_uid887
      port map ( clk  => clk,
                 X => tile_28_X,
                 Y => tile_28_Y,
                 R => tile_28_output);

tile_28_filtered_output <= tile_28_output(3 downto 0);
   bh793_w73_4 <= tile_28_filtered_output(0);
   bh793_w74_4 <= tile_28_filtered_output(1);
   bh793_w75_4 <= tile_28_filtered_output(2);
   bh793_w76_4 <= tile_28_filtered_output(3);
   tile_29_X <= X(20 downto 17);
   tile_29_Y <= Y(52 downto 52);
   tile_29_mult: IntMultiplierLUT_4x1_F200_uid889
      port map ( clk  => clk,
                 X => tile_29_X,
                 Y => tile_29_Y,
                 R => tile_29_output);

tile_29_filtered_output <= tile_29_output(3 downto 0);
   bh793_w69_4 <= tile_29_filtered_output(0);
   bh793_w70_4 <= tile_29_filtered_output(1);
   bh793_w71_4 <= tile_29_filtered_output(2);
   bh793_w72_4 <= tile_29_filtered_output(3);
   tile_30_X <= X(33 downto 32);
   tile_30_Y <= Y(51 downto 50);
   tile_30_mult: IntMultiplierLUT_2x2_F200_uid891
      port map ( clk  => clk,
                 X => tile_30_X,
                 Y => tile_30_Y,
                 R => tile_30_output);

tile_30_filtered_output <= tile_30_output(3 downto 0);
   bh793_w82_3 <= tile_30_filtered_output(0);
   bh793_w83_3 <= tile_30_filtered_output(1);
   bh793_w84_3 <= tile_30_filtered_output(2);
   bh793_w85_3 <= tile_30_filtered_output(3);
   tile_31_X <= X(31 downto 29);
   tile_31_Y <= Y(51 downto 50);
   tile_31_mult: IntMultiplierLUT_3x2_F200_uid896
      port map ( clk  => clk,
                 X => tile_31_X,
                 Y => tile_31_Y,
                 R => tile_31_output);

tile_31_filtered_output <= tile_31_output(4 downto 0);
   bh793_w79_4 <= tile_31_filtered_output(0);
   bh793_w80_4 <= tile_31_filtered_output(1);
   bh793_w81_4 <= tile_31_filtered_output(2);
   bh793_w82_4 <= tile_31_filtered_output(3);
   bh793_w83_4 <= tile_31_filtered_output(4);
   tile_32_X <= X(28 downto 26);
   tile_32_Y <= Y(51 downto 50);
   tile_32_mult: IntMultiplierLUT_3x2_F200_uid901
      port map ( clk  => clk,
                 X => tile_32_X,
                 Y => tile_32_Y,
                 R => tile_32_output);

tile_32_filtered_output <= tile_32_output(4 downto 0);
   bh793_w76_5 <= tile_32_filtered_output(0);
   bh793_w77_4 <= tile_32_filtered_output(1);
   bh793_w78_4 <= tile_32_filtered_output(2);
   bh793_w79_5 <= tile_32_filtered_output(3);
   bh793_w80_5 <= tile_32_filtered_output(4);
   tile_33_X <= X(25 downto 23);
   tile_33_Y <= Y(51 downto 50);
   tile_33_mult: IntMultiplierLUT_3x2_F200_uid906
      port map ( clk  => clk,
                 X => tile_33_X,
                 Y => tile_33_Y,
                 R => tile_33_output);

tile_33_filtered_output <= tile_33_output(4 downto 0);
   bh793_w73_5 <= tile_33_filtered_output(0);
   bh793_w74_5 <= tile_33_filtered_output(1);
   bh793_w75_5 <= tile_33_filtered_output(2);
   bh793_w76_6 <= tile_33_filtered_output(3);
   bh793_w77_5 <= tile_33_filtered_output(4);
   tile_34_X <= X(22 downto 20);
   tile_34_Y <= Y(51 downto 50);
   tile_34_mult: IntMultiplierLUT_3x2_F200_uid911
      port map ( clk  => clk,
                 X => tile_34_X,
                 Y => tile_34_Y,
                 R => tile_34_output);

tile_34_filtered_output <= tile_34_output(4 downto 0);
   bh793_w70_5 <= tile_34_filtered_output(0);
   bh793_w71_5 <= tile_34_filtered_output(1);
   bh793_w72_5 <= tile_34_filtered_output(2);
   bh793_w73_6 <= tile_34_filtered_output(3);
   bh793_w74_6 <= tile_34_filtered_output(4);
   tile_35_X <= X(19 downto 17);
   tile_35_Y <= Y(51 downto 50);
   tile_35_mult: IntMultiplierLUT_3x2_F200_uid916
      port map ( clk  => clk,
                 X => tile_35_X,
                 Y => tile_35_Y,
                 R => tile_35_output);

tile_35_filtered_output <= tile_35_output(4 downto 0);
   bh793_w67_6 <= tile_35_filtered_output(0);
   bh793_w68_6 <= tile_35_filtered_output(1);
   bh793_w69_5 <= tile_35_filtered_output(2);
   bh793_w70_6 <= tile_35_filtered_output(3);
   bh793_w71_6 <= tile_35_filtered_output(4);
   tile_36_X <= X(33 downto 32);
   tile_36_Y <= Y(49 downto 48);
   tile_36_mult: IntMultiplierLUT_2x2_F200_uid921
      port map ( clk  => clk,
                 X => tile_36_X,
                 Y => tile_36_Y,
                 R => tile_36_output);

tile_36_filtered_output <= tile_36_output(3 downto 0);
   bh793_w80_6 <= tile_36_filtered_output(0);
   bh793_w81_5 <= tile_36_filtered_output(1);
   bh793_w82_5 <= tile_36_filtered_output(2);
   bh793_w83_5 <= tile_36_filtered_output(3);
   tile_37_X <= X(31 downto 29);
   tile_37_Y <= Y(49 downto 48);
   tile_37_mult: IntMultiplierLUT_3x2_F200_uid926
      port map ( clk  => clk,
                 X => tile_37_X,
                 Y => tile_37_Y,
                 R => tile_37_output);

tile_37_filtered_output <= tile_37_output(4 downto 0);
   bh793_w77_6 <= tile_37_filtered_output(0);
   bh793_w78_5 <= tile_37_filtered_output(1);
   bh793_w79_6 <= tile_37_filtered_output(2);
   bh793_w80_7 <= tile_37_filtered_output(3);
   bh793_w81_6 <= tile_37_filtered_output(4);
   tile_38_X <= X(28 downto 26);
   tile_38_Y <= Y(49 downto 48);
   tile_38_mult: IntMultiplierLUT_3x2_F200_uid931
      port map ( clk  => clk,
                 X => tile_38_X,
                 Y => tile_38_Y,
                 R => tile_38_output);

tile_38_filtered_output <= tile_38_output(4 downto 0);
   bh793_w74_7 <= tile_38_filtered_output(0);
   bh793_w75_6 <= tile_38_filtered_output(1);
   bh793_w76_7 <= tile_38_filtered_output(2);
   bh793_w77_7 <= tile_38_filtered_output(3);
   bh793_w78_6 <= tile_38_filtered_output(4);
   tile_39_X <= X(25 downto 23);
   tile_39_Y <= Y(49 downto 48);
   tile_39_mult: IntMultiplierLUT_3x2_F200_uid936
      port map ( clk  => clk,
                 X => tile_39_X,
                 Y => tile_39_Y,
                 R => tile_39_output);

tile_39_filtered_output <= tile_39_output(4 downto 0);
   bh793_w71_7 <= tile_39_filtered_output(0);
   bh793_w72_6 <= tile_39_filtered_output(1);
   bh793_w73_7 <= tile_39_filtered_output(2);
   bh793_w74_8 <= tile_39_filtered_output(3);
   bh793_w75_7 <= tile_39_filtered_output(4);
   tile_40_X <= X(22 downto 20);
   tile_40_Y <= Y(49 downto 48);
   tile_40_mult: IntMultiplierLUT_3x2_F200_uid941
      port map ( clk  => clk,
                 X => tile_40_X,
                 Y => tile_40_Y,
                 R => tile_40_output);

tile_40_filtered_output <= tile_40_output(4 downto 0);
   bh793_w68_7 <= tile_40_filtered_output(0);
   bh793_w69_6 <= tile_40_filtered_output(1);
   bh793_w70_7 <= tile_40_filtered_output(2);
   bh793_w71_8 <= tile_40_filtered_output(3);
   bh793_w72_7 <= tile_40_filtered_output(4);
   tile_41_X <= X(19 downto 17);
   tile_41_Y <= Y(49 downto 48);
   tile_41_mult: IntMultiplierLUT_3x2_F200_uid946
      port map ( clk  => clk,
                 X => tile_41_X,
                 Y => tile_41_Y,
                 R => tile_41_output);

tile_41_filtered_output <= tile_41_output(4 downto 0);
   bh793_w65_8 <= tile_41_filtered_output(0);
   bh793_w66_8 <= tile_41_filtered_output(1);
   bh793_w67_7 <= tile_41_filtered_output(2);
   bh793_w68_8 <= tile_41_filtered_output(3);
   bh793_w69_7 <= tile_41_filtered_output(4);
   tile_42_X <= X(50 downto 50);
   tile_42_Y <= Y(52 downto 52);
   tile_42_mult: IntMultiplierLUT_1x1_F200_uid951
      port map ( clk  => clk,
                 X => tile_42_X,
                 Y => tile_42_Y,
                 R => tile_42_output);

tile_42_filtered_output <= tile_42_output(0 downto 0);
   bh793_w102_0 <= tile_42_filtered_output(0);
   tile_43_X <= X(49 downto 46);
   tile_43_Y <= Y(52 downto 52);
   tile_43_mult: IntMultiplierLUT_4x1_F200_uid953
      port map ( clk  => clk,
                 X => tile_43_X,
                 Y => tile_43_Y,
                 R => tile_43_output);

tile_43_filtered_output <= tile_43_output(3 downto 0);
   bh793_w98_2 <= tile_43_filtered_output(0);
   bh793_w99_1 <= tile_43_filtered_output(1);
   bh793_w100_1 <= tile_43_filtered_output(2);
   bh793_w101_0 <= tile_43_filtered_output(3);
   tile_44_X <= X(45 downto 42);
   tile_44_Y <= Y(52 downto 52);
   tile_44_mult: IntMultiplierLUT_4x1_F200_uid955
      port map ( clk  => clk,
                 X => tile_44_X,
                 Y => tile_44_Y,
                 R => tile_44_output);

tile_44_filtered_output <= tile_44_output(3 downto 0);
   bh793_w94_2 <= tile_44_filtered_output(0);
   bh793_w95_2 <= tile_44_filtered_output(1);
   bh793_w96_2 <= tile_44_filtered_output(2);
   bh793_w97_2 <= tile_44_filtered_output(3);
   tile_45_X <= X(41 downto 38);
   tile_45_Y <= Y(52 downto 52);
   tile_45_mult: IntMultiplierLUT_4x1_F200_uid957
      port map ( clk  => clk,
                 X => tile_45_X,
                 Y => tile_45_Y,
                 R => tile_45_output);

tile_45_filtered_output <= tile_45_output(3 downto 0);
   bh793_w90_2 <= tile_45_filtered_output(0);
   bh793_w91_2 <= tile_45_filtered_output(1);
   bh793_w92_2 <= tile_45_filtered_output(2);
   bh793_w93_2 <= tile_45_filtered_output(3);
   tile_46_X <= X(37 downto 34);
   tile_46_Y <= Y(52 downto 52);
   tile_46_mult: IntMultiplierLUT_4x1_F200_uid959
      port map ( clk  => clk,
                 X => tile_46_X,
                 Y => tile_46_Y,
                 R => tile_46_output);

tile_46_filtered_output <= tile_46_output(3 downto 0);
   bh793_w86_2 <= tile_46_filtered_output(0);
   bh793_w87_2 <= tile_46_filtered_output(1);
   bh793_w88_2 <= tile_46_filtered_output(2);
   bh793_w89_2 <= tile_46_filtered_output(3);
   tile_47_X <= X(50 downto 49);
   tile_47_Y <= Y(51 downto 50);
   tile_47_mult: IntMultiplierLUT_2x2_F200_uid961
      port map ( clk  => clk,
                 X => tile_47_X,
                 Y => tile_47_Y,
                 R => tile_47_output);

tile_47_filtered_output <= tile_47_output(3 downto 0);
   bh793_w99_2 <= tile_47_filtered_output(0);
   bh793_w100_2 <= tile_47_filtered_output(1);
   bh793_w101_1 <= tile_47_filtered_output(2);
   bh793_w102_1 <= tile_47_filtered_output(3);
   tile_48_X <= X(48 downto 46);
   tile_48_Y <= Y(51 downto 50);
   tile_48_mult: IntMultiplierLUT_3x2_F200_uid966
      port map ( clk  => clk,
                 X => tile_48_X,
                 Y => tile_48_Y,
                 R => tile_48_output);

tile_48_filtered_output <= tile_48_output(4 downto 0);
   bh793_w96_3 <= tile_48_filtered_output(0);
   bh793_w97_3 <= tile_48_filtered_output(1);
   bh793_w98_3 <= tile_48_filtered_output(2);
   bh793_w99_3 <= tile_48_filtered_output(3);
   bh793_w100_3 <= tile_48_filtered_output(4);
   tile_49_X <= X(45 downto 43);
   tile_49_Y <= Y(51 downto 50);
   tile_49_mult: IntMultiplierLUT_3x2_F200_uid971
      port map ( clk  => clk,
                 X => tile_49_X,
                 Y => tile_49_Y,
                 R => tile_49_output);

tile_49_filtered_output <= tile_49_output(4 downto 0);
   bh793_w93_3 <= tile_49_filtered_output(0);
   bh793_w94_3 <= tile_49_filtered_output(1);
   bh793_w95_3 <= tile_49_filtered_output(2);
   bh793_w96_4 <= tile_49_filtered_output(3);
   bh793_w97_4 <= tile_49_filtered_output(4);
   tile_50_X <= X(42 downto 40);
   tile_50_Y <= Y(51 downto 50);
   tile_50_mult: IntMultiplierLUT_3x2_F200_uid976
      port map ( clk  => clk,
                 X => tile_50_X,
                 Y => tile_50_Y,
                 R => tile_50_output);

tile_50_filtered_output <= tile_50_output(4 downto 0);
   bh793_w90_3 <= tile_50_filtered_output(0);
   bh793_w91_3 <= tile_50_filtered_output(1);
   bh793_w92_3 <= tile_50_filtered_output(2);
   bh793_w93_4 <= tile_50_filtered_output(3);
   bh793_w94_4 <= tile_50_filtered_output(4);
   tile_51_X <= X(39 downto 37);
   tile_51_Y <= Y(51 downto 50);
   tile_51_mult: IntMultiplierLUT_3x2_F200_uid981
      port map ( clk  => clk,
                 X => tile_51_X,
                 Y => tile_51_Y,
                 R => tile_51_output);

tile_51_filtered_output <= tile_51_output(4 downto 0);
   bh793_w87_3 <= tile_51_filtered_output(0);
   bh793_w88_3 <= tile_51_filtered_output(1);
   bh793_w89_3 <= tile_51_filtered_output(2);
   bh793_w90_4 <= tile_51_filtered_output(3);
   bh793_w91_4 <= tile_51_filtered_output(4);
   tile_52_X <= X(36 downto 34);
   tile_52_Y <= Y(51 downto 50);
   tile_52_mult: IntMultiplierLUT_3x2_F200_uid986
      port map ( clk  => clk,
                 X => tile_52_X,
                 Y => tile_52_Y,
                 R => tile_52_output);

tile_52_filtered_output <= tile_52_output(4 downto 0);
   bh793_w84_4 <= tile_52_filtered_output(0);
   bh793_w85_4 <= tile_52_filtered_output(1);
   bh793_w86_3 <= tile_52_filtered_output(2);
   bh793_w87_4 <= tile_52_filtered_output(3);
   bh793_w88_4 <= tile_52_filtered_output(4);
   tile_53_X <= X(50 downto 49);
   tile_53_Y <= Y(49 downto 48);
   tile_53_mult: IntMultiplierLUT_2x2_F200_uid991
      port map ( clk  => clk,
                 X => tile_53_X,
                 Y => tile_53_Y,
                 R => tile_53_output);

tile_53_filtered_output <= tile_53_output(3 downto 0);
   bh793_w97_5 <= tile_53_filtered_output(0);
   bh793_w98_4 <= tile_53_filtered_output(1);
   bh793_w99_4 <= tile_53_filtered_output(2);
   bh793_w100_4 <= tile_53_filtered_output(3);
   tile_54_X <= X(48 downto 46);
   tile_54_Y <= Y(49 downto 48);
   tile_54_mult: IntMultiplierLUT_3x2_F200_uid996
      port map ( clk  => clk,
                 X => tile_54_X,
                 Y => tile_54_Y,
                 R => tile_54_output);

tile_54_filtered_output <= tile_54_output(4 downto 0);
   bh793_w94_5 <= tile_54_filtered_output(0);
   bh793_w95_4 <= tile_54_filtered_output(1);
   bh793_w96_5 <= tile_54_filtered_output(2);
   bh793_w97_6 <= tile_54_filtered_output(3);
   bh793_w98_5 <= tile_54_filtered_output(4);
   tile_55_X <= X(45 downto 43);
   tile_55_Y <= Y(49 downto 48);
   tile_55_mult: IntMultiplierLUT_3x2_F200_uid1001
      port map ( clk  => clk,
                 X => tile_55_X,
                 Y => tile_55_Y,
                 R => tile_55_output);

tile_55_filtered_output <= tile_55_output(4 downto 0);
   bh793_w91_5 <= tile_55_filtered_output(0);
   bh793_w92_4 <= tile_55_filtered_output(1);
   bh793_w93_5 <= tile_55_filtered_output(2);
   bh793_w94_6 <= tile_55_filtered_output(3);
   bh793_w95_5 <= tile_55_filtered_output(4);
   tile_56_X <= X(42 downto 40);
   tile_56_Y <= Y(49 downto 48);
   tile_56_mult: IntMultiplierLUT_3x2_F200_uid1006
      port map ( clk  => clk,
                 X => tile_56_X,
                 Y => tile_56_Y,
                 R => tile_56_output);

tile_56_filtered_output <= tile_56_output(4 downto 0);
   bh793_w88_5 <= tile_56_filtered_output(0);
   bh793_w89_4 <= tile_56_filtered_output(1);
   bh793_w90_5 <= tile_56_filtered_output(2);
   bh793_w91_6 <= tile_56_filtered_output(3);
   bh793_w92_5 <= tile_56_filtered_output(4);
   tile_57_X <= X(39 downto 37);
   tile_57_Y <= Y(49 downto 48);
   tile_57_mult: IntMultiplierLUT_3x2_F200_uid1011
      port map ( clk  => clk,
                 X => tile_57_X,
                 Y => tile_57_Y,
                 R => tile_57_output);

tile_57_filtered_output <= tile_57_output(4 downto 0);
   bh793_w85_5 <= tile_57_filtered_output(0);
   bh793_w86_4 <= tile_57_filtered_output(1);
   bh793_w87_5 <= tile_57_filtered_output(2);
   bh793_w88_6 <= tile_57_filtered_output(3);
   bh793_w89_5 <= tile_57_filtered_output(4);
   tile_58_X <= X(36 downto 34);
   tile_58_Y <= Y(49 downto 48);
   tile_58_mult: IntMultiplierLUT_3x2_F200_uid1016
      port map ( clk  => clk,
                 X => tile_58_X,
                 Y => tile_58_Y,
                 R => tile_58_output);

tile_58_filtered_output <= tile_58_output(4 downto 0);
   bh793_w82_6 <= tile_58_filtered_output(0);
   bh793_w83_6 <= tile_58_filtered_output(1);
   bh793_w84_5 <= tile_58_filtered_output(2);
   bh793_w85_6 <= tile_58_filtered_output(3);
   bh793_w86_5 <= tile_58_filtered_output(4);
   tile_59_X <= X(52 downto 51);
   tile_59_Y <= Y(52 downto 51);
   tile_59_mult: IntMultiplierLUT_2x2_F200_uid1021
      port map ( clk  => clk,
                 X => tile_59_X,
                 Y => tile_59_Y,
                 R => tile_59_output);

tile_59_filtered_output <= tile_59_output(3 downto 0);
   bh793_w102_2 <= tile_59_filtered_output(0);
   bh793_w103_0 <= tile_59_filtered_output(1);
   bh793_w104_0 <= tile_59_filtered_output(2);
   bh793_w105_0 <= tile_59_filtered_output(3);
   tile_60_X <= X(52 downto 51);
   tile_60_Y <= Y(50 downto 48);
   tile_60_mult: IntMultiplierLUT_2x3_F200_uid1026
      port map ( clk  => clk,
                 X => tile_60_X,
                 Y => tile_60_Y,
                 R => tile_60_output);

tile_60_filtered_output <= tile_60_output(4 downto 0);
   bh793_w99_5 <= tile_60_filtered_output(0);
   bh793_w100_5 <= tile_60_filtered_output(1);
   bh793_w101_2 <= tile_60_filtered_output(2);
   bh793_w102_3 <= tile_60_filtered_output(3);
   bh793_w103_1 <= tile_60_filtered_output(4);

   -- Adding the constant bits
      -- All the constant bits are zero, nothing to add


   Compressor_23_3_F200_uid1032_bh793_uid1033_In0 <= "" & bh793_w17_0 & bh793_w17_1 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1033_In1 <= "" & bh793_w18_0 & bh793_w18_1;
   Compressor_23_3_F200_uid1032_uid1033: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1033_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1033_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1033_Out0_copy1034);
   Compressor_23_3_F200_uid1032_bh793_uid1033_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1033_Out0_copy1034; -- output copy to hold a pipeline register if needed

   bh793_w17_2 <= Compressor_23_3_F200_uid1032_bh793_uid1033_Out0(0);
   bh793_w18_2 <= Compressor_23_3_F200_uid1032_bh793_uid1033_Out0(1);
   bh793_w19_2 <= Compressor_23_3_F200_uid1032_bh793_uid1033_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1035_In0 <= "" & bh793_w19_0 & bh793_w19_1 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1035_In1 <= "" & bh793_w20_0 & bh793_w20_1;
   Compressor_23_3_F200_uid1032_uid1035: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1035_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1035_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1035_Out0_copy1036);
   Compressor_23_3_F200_uid1032_bh793_uid1035_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1035_Out0_copy1036; -- output copy to hold a pipeline register if needed

   bh793_w19_3 <= Compressor_23_3_F200_uid1032_bh793_uid1035_Out0(0);
   bh793_w20_2 <= Compressor_23_3_F200_uid1032_bh793_uid1035_Out0(1);
   bh793_w21_2 <= Compressor_23_3_F200_uid1032_bh793_uid1035_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1037_In0 <= "" & bh793_w21_0 & bh793_w21_1 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1037_In1 <= "" & bh793_w22_0 & bh793_w22_1;
   Compressor_23_3_F200_uid1032_uid1037: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1037_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1037_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1037_Out0_copy1038);
   Compressor_23_3_F200_uid1032_bh793_uid1037_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1037_Out0_copy1038; -- output copy to hold a pipeline register if needed

   bh793_w21_3 <= Compressor_23_3_F200_uid1032_bh793_uid1037_Out0(0);
   bh793_w22_2 <= Compressor_23_3_F200_uid1032_bh793_uid1037_Out0(1);
   bh793_w23_2 <= Compressor_23_3_F200_uid1032_bh793_uid1037_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1041_In0 <= "" & bh793_w23_0 & bh793_w23_1 & "0";
   Compressor_3_2_F200_uid1040_uid1041: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1041_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1041_Out0_copy1042);
   Compressor_3_2_F200_uid1040_bh793_uid1041_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1041_Out0_copy1042; -- output copy to hold a pipeline register if needed

   bh793_w23_3 <= Compressor_3_2_F200_uid1040_bh793_uid1041_Out0(0);
   bh793_w24_3 <= Compressor_3_2_F200_uid1040_bh793_uid1041_Out0(1);

   Compressor_23_3_F200_uid1032_bh793_uid1043_In0 <= "" & bh793_w24_0 & bh793_w24_1 & bh793_w24_2;
   Compressor_23_3_F200_uid1032_bh793_uid1043_In1 <= "" & bh793_w25_0 & bh793_w25_1;
   Compressor_23_3_F200_uid1032_uid1043: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1043_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1043_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1043_Out0_copy1044);
   Compressor_23_3_F200_uid1032_bh793_uid1043_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1043_Out0_copy1044; -- output copy to hold a pipeline register if needed

   bh793_w24_4 <= Compressor_23_3_F200_uid1032_bh793_uid1043_Out0(0);
   bh793_w25_3 <= Compressor_23_3_F200_uid1032_bh793_uid1043_Out0(1);
   bh793_w26_3 <= Compressor_23_3_F200_uid1032_bh793_uid1043_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1045_In0 <= "" & bh793_w26_0 & bh793_w26_1 & bh793_w26_2;
   Compressor_23_3_F200_uid1032_bh793_uid1045_In1 <= "" & bh793_w27_0 & bh793_w27_1;
   Compressor_23_3_F200_uid1032_uid1045: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1045_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1045_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1045_Out0_copy1046);
   Compressor_23_3_F200_uid1032_bh793_uid1045_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1045_Out0_copy1046; -- output copy to hold a pipeline register if needed

   bh793_w26_4 <= Compressor_23_3_F200_uid1032_bh793_uid1045_Out0(0);
   bh793_w27_3 <= Compressor_23_3_F200_uid1032_bh793_uid1045_Out0(1);
   bh793_w28_3 <= Compressor_23_3_F200_uid1032_bh793_uid1045_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1047_In0 <= "" & bh793_w28_0 & bh793_w28_1 & bh793_w28_2;
   Compressor_23_3_F200_uid1032_bh793_uid1047_In1 <= "" & bh793_w29_0 & bh793_w29_1;
   Compressor_23_3_F200_uid1032_uid1047: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1047_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1047_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1047_Out0_copy1048);
   Compressor_23_3_F200_uid1032_bh793_uid1047_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1047_Out0_copy1048; -- output copy to hold a pipeline register if needed

   bh793_w28_4 <= Compressor_23_3_F200_uid1032_bh793_uid1047_Out0(0);
   bh793_w29_3 <= Compressor_23_3_F200_uid1032_bh793_uid1047_Out0(1);
   bh793_w30_3 <= Compressor_23_3_F200_uid1032_bh793_uid1047_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1049_In0 <= "" & bh793_w30_0 & bh793_w30_1 & bh793_w30_2;
   Compressor_23_3_F200_uid1032_bh793_uid1049_In1 <= "" & bh793_w31_0 & bh793_w31_1;
   Compressor_23_3_F200_uid1032_uid1049: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1049_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1049_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1049_Out0_copy1050);
   Compressor_23_3_F200_uid1032_bh793_uid1049_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1049_Out0_copy1050; -- output copy to hold a pipeline register if needed

   bh793_w30_4 <= Compressor_23_3_F200_uid1032_bh793_uid1049_Out0(0);
   bh793_w31_3 <= Compressor_23_3_F200_uid1032_bh793_uid1049_Out0(1);
   bh793_w32_3 <= Compressor_23_3_F200_uid1032_bh793_uid1049_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1051_In0 <= "" & bh793_w32_0 & bh793_w32_1 & bh793_w32_2;
   Compressor_23_3_F200_uid1032_bh793_uid1051_In1 <= "" & bh793_w33_0 & bh793_w33_1;
   Compressor_23_3_F200_uid1032_uid1051: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1051_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1051_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1051_Out0_copy1052);
   Compressor_23_3_F200_uid1032_bh793_uid1051_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1051_Out0_copy1052; -- output copy to hold a pipeline register if needed

   bh793_w32_4 <= Compressor_23_3_F200_uid1032_bh793_uid1051_Out0(0);
   bh793_w33_3 <= Compressor_23_3_F200_uid1032_bh793_uid1051_Out0(1);
   bh793_w34_4 <= Compressor_23_3_F200_uid1032_bh793_uid1051_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1055_In0 <= "" & bh793_w34_0 & bh793_w34_1 & bh793_w34_2 & bh793_w34_3;
   Compressor_14_3_F200_uid1054_bh793_uid1055_In1 <= "" & bh793_w35_0;
   Compressor_14_3_F200_uid1054_uid1055: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1055_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1055_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1055_Out0_copy1056);
   Compressor_14_3_F200_uid1054_bh793_uid1055_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1055_Out0_copy1056; -- output copy to hold a pipeline register if needed

   bh793_w34_5 <= Compressor_14_3_F200_uid1054_bh793_uid1055_Out0(0);
   bh793_w35_4 <= Compressor_14_3_F200_uid1054_bh793_uid1055_Out0(1);
   bh793_w36_4 <= Compressor_14_3_F200_uid1054_bh793_uid1055_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1057_In0 <= "" & bh793_w35_1 & bh793_w35_2 & bh793_w35_3;
   Compressor_3_2_F200_uid1040_uid1057: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1057_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1057_Out0_copy1058);
   Compressor_3_2_F200_uid1040_bh793_uid1057_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1057_Out0_copy1058; -- output copy to hold a pipeline register if needed

   bh793_w35_5 <= Compressor_3_2_F200_uid1040_bh793_uid1057_Out0(0);
   bh793_w36_5 <= Compressor_3_2_F200_uid1040_bh793_uid1057_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1059_In0 <= "" & bh793_w36_0 & bh793_w36_1 & bh793_w36_2 & bh793_w36_3;
   Compressor_14_3_F200_uid1054_bh793_uid1059_In1 <= "" & bh793_w37_0;
   Compressor_14_3_F200_uid1054_uid1059: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1059_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1059_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1059_Out0_copy1060);
   Compressor_14_3_F200_uid1054_bh793_uid1059_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1059_Out0_copy1060; -- output copy to hold a pipeline register if needed

   bh793_w36_6 <= Compressor_14_3_F200_uid1054_bh793_uid1059_Out0(0);
   bh793_w37_4 <= Compressor_14_3_F200_uid1054_bh793_uid1059_Out0(1);
   bh793_w38_4 <= Compressor_14_3_F200_uid1054_bh793_uid1059_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1061_In0 <= "" & bh793_w37_1 & bh793_w37_2 & bh793_w37_3;
   Compressor_3_2_F200_uid1040_uid1061: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1061_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1061_Out0_copy1062);
   Compressor_3_2_F200_uid1040_bh793_uid1061_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1061_Out0_copy1062; -- output copy to hold a pipeline register if needed

   bh793_w37_5 <= Compressor_3_2_F200_uid1040_bh793_uid1061_Out0(0);
   bh793_w38_5 <= Compressor_3_2_F200_uid1040_bh793_uid1061_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1063_In0 <= "" & bh793_w38_0 & bh793_w38_1 & bh793_w38_2 & bh793_w38_3;
   Compressor_14_3_F200_uid1054_bh793_uid1063_In1 <= "" & bh793_w39_0;
   Compressor_14_3_F200_uid1054_uid1063: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1063_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1063_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1063_Out0_copy1064);
   Compressor_14_3_F200_uid1054_bh793_uid1063_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1063_Out0_copy1064; -- output copy to hold a pipeline register if needed

   bh793_w38_6 <= Compressor_14_3_F200_uid1054_bh793_uid1063_Out0(0);
   bh793_w39_4 <= Compressor_14_3_F200_uid1054_bh793_uid1063_Out0(1);
   bh793_w40_4 <= Compressor_14_3_F200_uid1054_bh793_uid1063_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1065_In0 <= "" & bh793_w39_1 & bh793_w39_2 & bh793_w39_3;
   Compressor_3_2_F200_uid1040_uid1065: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1065_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1065_Out0_copy1066);
   Compressor_3_2_F200_uid1040_bh793_uid1065_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1065_Out0_copy1066; -- output copy to hold a pipeline register if needed

   bh793_w39_5 <= Compressor_3_2_F200_uid1040_bh793_uid1065_Out0(0);
   bh793_w40_5 <= Compressor_3_2_F200_uid1040_bh793_uid1065_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1067_In0 <= "" & bh793_w40_0 & bh793_w40_1 & bh793_w40_2 & bh793_w40_3;
   Compressor_14_3_F200_uid1054_bh793_uid1067_In1 <= "" & bh793_w41_0;
   Compressor_14_3_F200_uid1054_uid1067: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1067_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1067_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1067_Out0_copy1068);
   Compressor_14_3_F200_uid1054_bh793_uid1067_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1067_Out0_copy1068; -- output copy to hold a pipeline register if needed

   bh793_w40_6 <= Compressor_14_3_F200_uid1054_bh793_uid1067_Out0(0);
   bh793_w41_4 <= Compressor_14_3_F200_uid1054_bh793_uid1067_Out0(1);
   bh793_w42_4 <= Compressor_14_3_F200_uid1054_bh793_uid1067_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1069_In0 <= "" & bh793_w41_1 & bh793_w41_2 & bh793_w41_3;
   Compressor_3_2_F200_uid1040_uid1069: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1069_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1069_Out0_copy1070);
   Compressor_3_2_F200_uid1040_bh793_uid1069_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1069_Out0_copy1070; -- output copy to hold a pipeline register if needed

   bh793_w41_5 <= Compressor_3_2_F200_uid1040_bh793_uid1069_Out0(0);
   bh793_w42_5 <= Compressor_3_2_F200_uid1040_bh793_uid1069_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1071_In0 <= "" & bh793_w42_0 & bh793_w42_1 & bh793_w42_2 & bh793_w42_3;
   Compressor_14_3_F200_uid1054_bh793_uid1071_In1 <= "" & bh793_w43_0;
   Compressor_14_3_F200_uid1054_uid1071: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1071_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1071_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1071_Out0_copy1072);
   Compressor_14_3_F200_uid1054_bh793_uid1071_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1071_Out0_copy1072; -- output copy to hold a pipeline register if needed

   bh793_w42_6 <= Compressor_14_3_F200_uid1054_bh793_uid1071_Out0(0);
   bh793_w43_4 <= Compressor_14_3_F200_uid1054_bh793_uid1071_Out0(1);
   bh793_w44_4 <= Compressor_14_3_F200_uid1054_bh793_uid1071_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1073_In0 <= "" & bh793_w43_1 & bh793_w43_2 & bh793_w43_3;
   Compressor_3_2_F200_uid1040_uid1073: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1073_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1073_Out0_copy1074);
   Compressor_3_2_F200_uid1040_bh793_uid1073_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1073_Out0_copy1074; -- output copy to hold a pipeline register if needed

   bh793_w43_5 <= Compressor_3_2_F200_uid1040_bh793_uid1073_Out0(0);
   bh793_w44_5 <= Compressor_3_2_F200_uid1040_bh793_uid1073_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1075_In0 <= "" & bh793_w44_0 & bh793_w44_1 & bh793_w44_2 & bh793_w44_3;
   Compressor_14_3_F200_uid1054_bh793_uid1075_In1 <= "" & bh793_w45_0;
   Compressor_14_3_F200_uid1054_uid1075: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1075_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1075_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1075_Out0_copy1076);
   Compressor_14_3_F200_uid1054_bh793_uid1075_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1075_Out0_copy1076; -- output copy to hold a pipeline register if needed

   bh793_w44_6 <= Compressor_14_3_F200_uid1054_bh793_uid1075_Out0(0);
   bh793_w45_4 <= Compressor_14_3_F200_uid1054_bh793_uid1075_Out0(1);
   bh793_w46_4 <= Compressor_14_3_F200_uid1054_bh793_uid1075_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1077_In0 <= "" & bh793_w45_1 & bh793_w45_2 & bh793_w45_3;
   Compressor_3_2_F200_uid1040_uid1077: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1077_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1077_Out0_copy1078);
   Compressor_3_2_F200_uid1040_bh793_uid1077_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1077_Out0_copy1078; -- output copy to hold a pipeline register if needed

   bh793_w45_5 <= Compressor_3_2_F200_uid1040_bh793_uid1077_Out0(0);
   bh793_w46_5 <= Compressor_3_2_F200_uid1040_bh793_uid1077_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1079_In0 <= "" & bh793_w46_0 & bh793_w46_1 & bh793_w46_2 & bh793_w46_3;
   Compressor_14_3_F200_uid1054_bh793_uid1079_In1 <= "" & bh793_w47_0;
   Compressor_14_3_F200_uid1054_uid1079: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1079_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1079_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1079_Out0_copy1080);
   Compressor_14_3_F200_uid1054_bh793_uid1079_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1079_Out0_copy1080; -- output copy to hold a pipeline register if needed

   bh793_w46_6 <= Compressor_14_3_F200_uid1054_bh793_uid1079_Out0(0);
   bh793_w47_4 <= Compressor_14_3_F200_uid1054_bh793_uid1079_Out0(1);
   bh793_w48_5 <= Compressor_14_3_F200_uid1054_bh793_uid1079_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1081_In0 <= "" & bh793_w47_1 & bh793_w47_2 & bh793_w47_3;
   Compressor_3_2_F200_uid1040_uid1081: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1081_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1081_Out0_copy1082);
   Compressor_3_2_F200_uid1040_bh793_uid1081_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1081_Out0_copy1082; -- output copy to hold a pipeline register if needed

   bh793_w47_5 <= Compressor_3_2_F200_uid1040_bh793_uid1081_Out0(0);
   bh793_w48_6 <= Compressor_3_2_F200_uid1040_bh793_uid1081_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1083_In0 <= "" & bh793_w48_0 & bh793_w48_1 & bh793_w48_2 & bh793_w48_3;
   Compressor_14_3_F200_uid1054_bh793_uid1083_In1 <= "" & bh793_w49_0;
   Compressor_14_3_F200_uid1054_uid1083: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1083_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1083_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1083_Out0_copy1084);
   Compressor_14_3_F200_uid1054_bh793_uid1083_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1083_Out0_copy1084; -- output copy to hold a pipeline register if needed

   bh793_w48_7 <= Compressor_14_3_F200_uid1054_bh793_uid1083_Out0(0);
   bh793_w49_5 <= Compressor_14_3_F200_uid1054_bh793_uid1083_Out0(1);
   bh793_w50_6 <= Compressor_14_3_F200_uid1054_bh793_uid1083_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1085_In0 <= "" & bh793_w49_1 & bh793_w49_2 & bh793_w49_3;
   Compressor_3_2_F200_uid1040_uid1085: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1085_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1085_Out0_copy1086);
   Compressor_3_2_F200_uid1040_bh793_uid1085_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1085_Out0_copy1086; -- output copy to hold a pipeline register if needed

   bh793_w49_6 <= Compressor_3_2_F200_uid1040_bh793_uid1085_Out0(0);
   bh793_w50_7 <= Compressor_3_2_F200_uid1040_bh793_uid1085_Out0(1);

   Compressor_6_3_F200_uid1088_bh793_uid1089_In0 <= "" & bh793_w50_0 & bh793_w50_1 & bh793_w50_2 & bh793_w50_3 & bh793_w50_4 & bh793_w50_5;
   Compressor_6_3_F200_uid1088_uid1089: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1089_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1089_Out0_copy1090);
   Compressor_6_3_F200_uid1088_bh793_uid1089_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1089_Out0_copy1090; -- output copy to hold a pipeline register if needed

   bh793_w50_8 <= Compressor_6_3_F200_uid1088_bh793_uid1089_Out0(0);
   bh793_w51_8 <= Compressor_6_3_F200_uid1088_bh793_uid1089_Out0(1);
   bh793_w52_9 <= Compressor_6_3_F200_uid1088_bh793_uid1089_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1091_In0 <= "" & bh793_w51_0 & bh793_w51_1 & bh793_w51_2 & bh793_w51_3 & bh793_w51_4 & "0";
   Compressor_6_3_F200_uid1088_uid1091: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1091_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1091_Out0_copy1092);
   Compressor_6_3_F200_uid1088_bh793_uid1091_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1091_Out0_copy1092; -- output copy to hold a pipeline register if needed

   bh793_w51_9 <= Compressor_6_3_F200_uid1088_bh793_uid1091_Out0(0);
   bh793_w52_10 <= Compressor_6_3_F200_uid1088_bh793_uid1091_Out0(1);
   bh793_w53_9 <= Compressor_6_3_F200_uid1088_bh793_uid1091_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1093_In0 <= "" & bh793_w51_5 & bh793_w51_6 & bh793_w51_7;
   Compressor_3_2_F200_uid1040_uid1093: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1093_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1093_Out0_copy1094);
   Compressor_3_2_F200_uid1040_bh793_uid1093_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1093_Out0_copy1094; -- output copy to hold a pipeline register if needed

   bh793_w51_10 <= Compressor_3_2_F200_uid1040_bh793_uid1093_Out0(0);
   bh793_w52_11 <= Compressor_3_2_F200_uid1040_bh793_uid1093_Out0(1);

   Compressor_6_3_F200_uid1088_bh793_uid1095_In0 <= "" & bh793_w52_0 & bh793_w52_1 & bh793_w52_2 & bh793_w52_3 & bh793_w52_4 & bh793_w52_5;
   Compressor_6_3_F200_uid1088_uid1095: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1095_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1095_Out0_copy1096);
   Compressor_6_3_F200_uid1088_bh793_uid1095_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1095_Out0_copy1096; -- output copy to hold a pipeline register if needed

   bh793_w52_12 <= Compressor_6_3_F200_uid1088_bh793_uid1095_Out0(0);
   bh793_w53_10 <= Compressor_6_3_F200_uid1088_bh793_uid1095_Out0(1);
   bh793_w54_10 <= Compressor_6_3_F200_uid1088_bh793_uid1095_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1097_In0 <= "" & bh793_w52_6 & bh793_w52_7 & bh793_w52_8;
   Compressor_23_3_F200_uid1032_bh793_uid1097_In1 <= "" & bh793_w53_0 & bh793_w53_1;
   Compressor_23_3_F200_uid1032_uid1097: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1097_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1097_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1097_Out0_copy1098);
   Compressor_23_3_F200_uid1032_bh793_uid1097_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1097_Out0_copy1098; -- output copy to hold a pipeline register if needed

   bh793_w52_13 <= Compressor_23_3_F200_uid1032_bh793_uid1097_Out0(0);
   bh793_w53_11 <= Compressor_23_3_F200_uid1032_bh793_uid1097_Out0(1);
   bh793_w54_11 <= Compressor_23_3_F200_uid1032_bh793_uid1097_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1099_In0 <= "" & bh793_w53_2 & bh793_w53_3 & bh793_w53_4 & bh793_w53_5 & bh793_w53_6 & bh793_w53_7;
   Compressor_6_3_F200_uid1088_uid1099: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1099_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1099_Out0_copy1100);
   Compressor_6_3_F200_uid1088_bh793_uid1099_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1099_Out0_copy1100; -- output copy to hold a pipeline register if needed

   bh793_w53_12 <= Compressor_6_3_F200_uid1088_bh793_uid1099_Out0(0);
   bh793_w54_12 <= Compressor_6_3_F200_uid1088_bh793_uid1099_Out0(1);
   bh793_w55_9 <= Compressor_6_3_F200_uid1088_bh793_uid1099_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1101_In0 <= "" & bh793_w54_0 & bh793_w54_1 & bh793_w54_2 & bh793_w54_3 & bh793_w54_4 & bh793_w54_5;
   Compressor_6_3_F200_uid1088_uid1101: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1101_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1101_Out0_copy1102);
   Compressor_6_3_F200_uid1088_bh793_uid1101_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1101_Out0_copy1102; -- output copy to hold a pipeline register if needed

   bh793_w54_13 <= Compressor_6_3_F200_uid1088_bh793_uid1101_Out0(0);
   bh793_w55_10 <= Compressor_6_3_F200_uid1088_bh793_uid1101_Out0(1);
   bh793_w56_9 <= Compressor_6_3_F200_uid1088_bh793_uid1101_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1103_In0 <= "" & bh793_w54_6 & bh793_w54_7 & bh793_w54_8 & bh793_w54_9;
   Compressor_14_3_F200_uid1054_bh793_uid1103_In1 <= "" & "0";
   Compressor_14_3_F200_uid1054_uid1103: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1103_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1103_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1103_Out0_copy1104);
   Compressor_14_3_F200_uid1054_bh793_uid1103_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1103_Out0_copy1104; -- output copy to hold a pipeline register if needed

   bh793_w54_14 <= Compressor_14_3_F200_uid1054_bh793_uid1103_Out0(0);
   bh793_w55_11 <= Compressor_14_3_F200_uid1054_bh793_uid1103_Out0(1);
   bh793_w56_10 <= Compressor_14_3_F200_uid1054_bh793_uid1103_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1105_In0 <= "" & bh793_w55_0 & bh793_w55_1 & bh793_w55_2 & bh793_w55_3 & bh793_w55_4 & bh793_w55_5;
   Compressor_6_3_F200_uid1088_uid1105: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1105_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1105_Out0_copy1106);
   Compressor_6_3_F200_uid1088_bh793_uid1105_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1105_Out0_copy1106; -- output copy to hold a pipeline register if needed

   bh793_w55_12 <= Compressor_6_3_F200_uid1088_bh793_uid1105_Out0(0);
   bh793_w56_11 <= Compressor_6_3_F200_uid1088_bh793_uid1105_Out0(1);
   bh793_w57_10 <= Compressor_6_3_F200_uid1088_bh793_uid1105_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1107_In0 <= "" & bh793_w55_6 & bh793_w55_7 & bh793_w55_8;
   Compressor_3_2_F200_uid1040_uid1107: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1107_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1107_Out0_copy1108);
   Compressor_3_2_F200_uid1040_bh793_uid1107_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1107_Out0_copy1108; -- output copy to hold a pipeline register if needed

   bh793_w55_13 <= Compressor_3_2_F200_uid1040_bh793_uid1107_Out0(0);
   bh793_w56_12 <= Compressor_3_2_F200_uid1040_bh793_uid1107_Out0(1);

   Compressor_6_3_F200_uid1088_bh793_uid1109_In0 <= "" & bh793_w56_0 & bh793_w56_1 & bh793_w56_2 & bh793_w56_3 & bh793_w56_4 & bh793_w56_5;
   Compressor_6_3_F200_uid1088_uid1109: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1109_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1109_Out0_copy1110);
   Compressor_6_3_F200_uid1088_bh793_uid1109_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1109_Out0_copy1110; -- output copy to hold a pipeline register if needed

   bh793_w56_13 <= Compressor_6_3_F200_uid1088_bh793_uid1109_Out0(0);
   bh793_w57_11 <= Compressor_6_3_F200_uid1088_bh793_uid1109_Out0(1);
   bh793_w58_9 <= Compressor_6_3_F200_uid1088_bh793_uid1109_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1111_In0 <= "" & bh793_w56_6 & bh793_w56_7 & bh793_w56_8;
   Compressor_3_2_F200_uid1040_uid1111: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1111_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1111_Out0_copy1112);
   Compressor_3_2_F200_uid1040_bh793_uid1111_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1111_Out0_copy1112; -- output copy to hold a pipeline register if needed

   bh793_w56_14 <= Compressor_3_2_F200_uid1040_bh793_uid1111_Out0(0);
   bh793_w57_12 <= Compressor_3_2_F200_uid1040_bh793_uid1111_Out0(1);

   Compressor_6_3_F200_uid1088_bh793_uid1113_In0 <= "" & bh793_w57_0 & bh793_w57_1 & bh793_w57_2 & bh793_w57_3 & bh793_w57_4 & bh793_w57_5;
   Compressor_6_3_F200_uid1088_uid1113: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1113_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1113_Out0_copy1114);
   Compressor_6_3_F200_uid1088_bh793_uid1113_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1113_Out0_copy1114; -- output copy to hold a pipeline register if needed

   bh793_w57_13 <= Compressor_6_3_F200_uid1088_bh793_uid1113_Out0(0);
   bh793_w58_10 <= Compressor_6_3_F200_uid1088_bh793_uid1113_Out0(1);
   bh793_w59_9 <= Compressor_6_3_F200_uid1088_bh793_uid1113_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1115_In0 <= "" & bh793_w57_6 & bh793_w57_7 & bh793_w57_8 & bh793_w57_9;
   Compressor_14_3_F200_uid1054_bh793_uid1115_In1 <= "" & "0";
   Compressor_14_3_F200_uid1054_uid1115: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1115_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1115_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1115_Out0_copy1116);
   Compressor_14_3_F200_uid1054_bh793_uid1115_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1115_Out0_copy1116; -- output copy to hold a pipeline register if needed

   bh793_w57_14 <= Compressor_14_3_F200_uid1054_bh793_uid1115_Out0(0);
   bh793_w58_11 <= Compressor_14_3_F200_uid1054_bh793_uid1115_Out0(1);
   bh793_w59_10 <= Compressor_14_3_F200_uid1054_bh793_uid1115_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1117_In0 <= "" & bh793_w58_0 & bh793_w58_1 & bh793_w58_2 & bh793_w58_3 & bh793_w58_4 & bh793_w58_5;
   Compressor_6_3_F200_uid1088_uid1117: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1117_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1117_Out0_copy1118);
   Compressor_6_3_F200_uid1088_bh793_uid1117_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1117_Out0_copy1118; -- output copy to hold a pipeline register if needed

   bh793_w58_12 <= Compressor_6_3_F200_uid1088_bh793_uid1117_Out0(0);
   bh793_w59_11 <= Compressor_6_3_F200_uid1088_bh793_uid1117_Out0(1);
   bh793_w60_10 <= Compressor_6_3_F200_uid1088_bh793_uid1117_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1119_In0 <= "" & bh793_w58_6 & bh793_w58_7 & bh793_w58_8;
   Compressor_3_2_F200_uid1040_uid1119: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1119_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1119_Out0_copy1120);
   Compressor_3_2_F200_uid1040_bh793_uid1119_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1119_Out0_copy1120; -- output copy to hold a pipeline register if needed

   bh793_w58_13 <= Compressor_3_2_F200_uid1040_bh793_uid1119_Out0(0);
   bh793_w59_12 <= Compressor_3_2_F200_uid1040_bh793_uid1119_Out0(1);

   Compressor_6_3_F200_uid1088_bh793_uid1121_In0 <= "" & bh793_w59_0 & bh793_w59_1 & bh793_w59_2 & bh793_w59_3 & bh793_w59_4 & bh793_w59_5;
   Compressor_6_3_F200_uid1088_uid1121: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1121_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1121_Out0_copy1122);
   Compressor_6_3_F200_uid1088_bh793_uid1121_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1121_Out0_copy1122; -- output copy to hold a pipeline register if needed

   bh793_w59_13 <= Compressor_6_3_F200_uid1088_bh793_uid1121_Out0(0);
   bh793_w60_11 <= Compressor_6_3_F200_uid1088_bh793_uid1121_Out0(1);
   bh793_w61_9 <= Compressor_6_3_F200_uid1088_bh793_uid1121_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1123_In0 <= "" & bh793_w59_6 & bh793_w59_7 & bh793_w59_8;
   Compressor_3_2_F200_uid1040_uid1123: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1123_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1123_Out0_copy1124);
   Compressor_3_2_F200_uid1040_bh793_uid1123_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1123_Out0_copy1124; -- output copy to hold a pipeline register if needed

   bh793_w59_14 <= Compressor_3_2_F200_uid1040_bh793_uid1123_Out0(0);
   bh793_w60_12 <= Compressor_3_2_F200_uid1040_bh793_uid1123_Out0(1);

   Compressor_6_3_F200_uid1088_bh793_uid1125_In0 <= "" & bh793_w60_0 & bh793_w60_1 & bh793_w60_2 & bh793_w60_3 & bh793_w60_4 & bh793_w60_5;
   Compressor_6_3_F200_uid1088_uid1125: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1125_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1125_Out0_copy1126);
   Compressor_6_3_F200_uid1088_bh793_uid1125_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1125_Out0_copy1126; -- output copy to hold a pipeline register if needed

   bh793_w60_13 <= Compressor_6_3_F200_uid1088_bh793_uid1125_Out0(0);
   bh793_w61_10 <= Compressor_6_3_F200_uid1088_bh793_uid1125_Out0(1);
   bh793_w62_9 <= Compressor_6_3_F200_uid1088_bh793_uid1125_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1127_In0 <= "" & bh793_w60_6 & bh793_w60_7 & bh793_w60_8 & bh793_w60_9;
   Compressor_14_3_F200_uid1054_bh793_uid1127_In1 <= "" & "0";
   Compressor_14_3_F200_uid1054_uid1127: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1127_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1127_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1127_Out0_copy1128);
   Compressor_14_3_F200_uid1054_bh793_uid1127_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1127_Out0_copy1128; -- output copy to hold a pipeline register if needed

   bh793_w60_14 <= Compressor_14_3_F200_uid1054_bh793_uid1127_Out0(0);
   bh793_w61_11 <= Compressor_14_3_F200_uid1054_bh793_uid1127_Out0(1);
   bh793_w62_10 <= Compressor_14_3_F200_uid1054_bh793_uid1127_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1129_In0 <= "" & bh793_w61_0 & bh793_w61_1 & bh793_w61_2 & bh793_w61_3 & bh793_w61_4 & bh793_w61_5;
   Compressor_6_3_F200_uid1088_uid1129: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1129_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1129_Out0_copy1130);
   Compressor_6_3_F200_uid1088_bh793_uid1129_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1129_Out0_copy1130; -- output copy to hold a pipeline register if needed

   bh793_w61_12 <= Compressor_6_3_F200_uid1088_bh793_uid1129_Out0(0);
   bh793_w62_11 <= Compressor_6_3_F200_uid1088_bh793_uid1129_Out0(1);
   bh793_w63_10 <= Compressor_6_3_F200_uid1088_bh793_uid1129_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1131_In0 <= "" & bh793_w61_6 & bh793_w61_7 & bh793_w61_8;
   Compressor_3_2_F200_uid1040_uid1131: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1131_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1131_Out0_copy1132);
   Compressor_3_2_F200_uid1040_bh793_uid1131_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1131_Out0_copy1132; -- output copy to hold a pipeline register if needed

   bh793_w61_13 <= Compressor_3_2_F200_uid1040_bh793_uid1131_Out0(0);
   bh793_w62_12 <= Compressor_3_2_F200_uid1040_bh793_uid1131_Out0(1);

   Compressor_6_3_F200_uid1088_bh793_uid1133_In0 <= "" & bh793_w62_0 & bh793_w62_1 & bh793_w62_2 & bh793_w62_3 & bh793_w62_4 & bh793_w62_5;
   Compressor_6_3_F200_uid1088_uid1133: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1133_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1133_Out0_copy1134);
   Compressor_6_3_F200_uid1088_bh793_uid1133_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1133_Out0_copy1134; -- output copy to hold a pipeline register if needed

   bh793_w62_13 <= Compressor_6_3_F200_uid1088_bh793_uid1133_Out0(0);
   bh793_w63_11 <= Compressor_6_3_F200_uid1088_bh793_uid1133_Out0(1);
   bh793_w64_9 <= Compressor_6_3_F200_uid1088_bh793_uid1133_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1135_In0 <= "" & bh793_w62_6 & bh793_w62_7 & bh793_w62_8;
   Compressor_3_2_F200_uid1040_uid1135: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1135_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1135_Out0_copy1136);
   Compressor_3_2_F200_uid1040_bh793_uid1135_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1135_Out0_copy1136; -- output copy to hold a pipeline register if needed

   bh793_w62_14 <= Compressor_3_2_F200_uid1040_bh793_uid1135_Out0(0);
   bh793_w63_12 <= Compressor_3_2_F200_uid1040_bh793_uid1135_Out0(1);

   Compressor_6_3_F200_uid1088_bh793_uid1137_In0 <= "" & bh793_w63_0 & bh793_w63_1 & bh793_w63_2 & bh793_w63_3 & bh793_w63_4 & bh793_w63_5;
   Compressor_6_3_F200_uid1088_uid1137: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1137_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1137_Out0_copy1138);
   Compressor_6_3_F200_uid1088_bh793_uid1137_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1137_Out0_copy1138; -- output copy to hold a pipeline register if needed

   bh793_w63_13 <= Compressor_6_3_F200_uid1088_bh793_uid1137_Out0(0);
   bh793_w64_10 <= Compressor_6_3_F200_uid1088_bh793_uid1137_Out0(1);
   bh793_w65_9 <= Compressor_6_3_F200_uid1088_bh793_uid1137_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1139_In0 <= "" & bh793_w63_6 & bh793_w63_7 & bh793_w63_8 & bh793_w63_9;
   Compressor_14_3_F200_uid1054_bh793_uid1139_In1 <= "" & "0";
   Compressor_14_3_F200_uid1054_uid1139: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1139_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1139_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1139_Out0_copy1140);
   Compressor_14_3_F200_uid1054_bh793_uid1139_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1139_Out0_copy1140; -- output copy to hold a pipeline register if needed

   bh793_w63_14 <= Compressor_14_3_F200_uid1054_bh793_uid1139_Out0(0);
   bh793_w64_11 <= Compressor_14_3_F200_uid1054_bh793_uid1139_Out0(1);
   bh793_w65_10 <= Compressor_14_3_F200_uid1054_bh793_uid1139_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1141_In0 <= "" & bh793_w64_0 & bh793_w64_1 & bh793_w64_2 & bh793_w64_3 & bh793_w64_4 & bh793_w64_5;
   Compressor_6_3_F200_uid1088_uid1141: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1141_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1141_Out0_copy1142);
   Compressor_6_3_F200_uid1088_bh793_uid1141_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1141_Out0_copy1142; -- output copy to hold a pipeline register if needed

   bh793_w64_12 <= Compressor_6_3_F200_uid1088_bh793_uid1141_Out0(0);
   bh793_w65_11 <= Compressor_6_3_F200_uid1088_bh793_uid1141_Out0(1);
   bh793_w66_9 <= Compressor_6_3_F200_uid1088_bh793_uid1141_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1143_In0 <= "" & bh793_w64_6 & bh793_w64_7 & bh793_w64_8;
   Compressor_3_2_F200_uid1040_uid1143: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1143_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1143_Out0_copy1144);
   Compressor_3_2_F200_uid1040_bh793_uid1143_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1143_Out0_copy1144; -- output copy to hold a pipeline register if needed

   bh793_w64_13 <= Compressor_3_2_F200_uid1040_bh793_uid1143_Out0(0);
   bh793_w65_12 <= Compressor_3_2_F200_uid1040_bh793_uid1143_Out0(1);

   Compressor_6_3_F200_uid1088_bh793_uid1145_In0 <= "" & bh793_w65_0 & bh793_w65_1 & bh793_w65_2 & bh793_w65_3 & bh793_w65_4 & bh793_w65_5;
   Compressor_6_3_F200_uid1088_uid1145: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1145_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1145_Out0_copy1146);
   Compressor_6_3_F200_uid1088_bh793_uid1145_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1145_Out0_copy1146; -- output copy to hold a pipeline register if needed

   bh793_w65_13 <= Compressor_6_3_F200_uid1088_bh793_uid1145_Out0(0);
   bh793_w66_10 <= Compressor_6_3_F200_uid1088_bh793_uid1145_Out0(1);
   bh793_w67_8 <= Compressor_6_3_F200_uid1088_bh793_uid1145_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1147_In0 <= "" & bh793_w65_6 & bh793_w65_7 & bh793_w65_8;
   Compressor_23_3_F200_uid1032_bh793_uid1147_In1 <= "" & "0" & "0";
   Compressor_23_3_F200_uid1032_uid1147: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1147_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1147_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1147_Out0_copy1148);
   Compressor_23_3_F200_uid1032_bh793_uid1147_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1147_Out0_copy1148; -- output copy to hold a pipeline register if needed

   bh793_w65_14 <= Compressor_23_3_F200_uid1032_bh793_uid1147_Out0(0);
   bh793_w66_11 <= Compressor_23_3_F200_uid1032_bh793_uid1147_Out0(1);
   bh793_w67_9 <= Compressor_23_3_F200_uid1032_bh793_uid1147_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1149_In0 <= "" & bh793_w66_0 & bh793_w66_1 & bh793_w66_2 & bh793_w66_3 & bh793_w66_4 & bh793_w66_5;
   Compressor_6_3_F200_uid1088_uid1149: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1149_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1149_Out0_copy1150);
   Compressor_6_3_F200_uid1088_bh793_uid1149_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1149_Out0_copy1150; -- output copy to hold a pipeline register if needed

   bh793_w66_12 <= Compressor_6_3_F200_uid1088_bh793_uid1149_Out0(0);
   bh793_w67_10 <= Compressor_6_3_F200_uid1088_bh793_uid1149_Out0(1);
   bh793_w68_9 <= Compressor_6_3_F200_uid1088_bh793_uid1149_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1151_In0 <= "" & bh793_w66_6 & bh793_w66_7 & bh793_w66_8;
   Compressor_23_3_F200_uid1032_bh793_uid1151_In1 <= "" & bh793_w67_0 & bh793_w67_1;
   Compressor_23_3_F200_uid1032_uid1151: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1151_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1151_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1151_Out0_copy1152);
   Compressor_23_3_F200_uid1032_bh793_uid1151_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1151_Out0_copy1152; -- output copy to hold a pipeline register if needed

   bh793_w66_13 <= Compressor_23_3_F200_uid1032_bh793_uid1151_Out0(0);
   bh793_w67_11 <= Compressor_23_3_F200_uid1032_bh793_uid1151_Out0(1);
   bh793_w68_10 <= Compressor_23_3_F200_uid1032_bh793_uid1151_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1153_In0 <= "" & bh793_w67_2 & bh793_w67_3 & bh793_w67_4 & bh793_w67_5 & bh793_w67_6 & bh793_w67_7;
   Compressor_6_3_F200_uid1088_uid1153: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1153_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1153_Out0_copy1154);
   Compressor_6_3_F200_uid1088_bh793_uid1153_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1153_Out0_copy1154; -- output copy to hold a pipeline register if needed

   bh793_w67_12 <= Compressor_6_3_F200_uid1088_bh793_uid1153_Out0(0);
   bh793_w68_11 <= Compressor_6_3_F200_uid1088_bh793_uid1153_Out0(1);
   bh793_w69_8 <= Compressor_6_3_F200_uid1088_bh793_uid1153_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1155_In0 <= "" & bh793_w68_0 & bh793_w68_1 & bh793_w68_2 & bh793_w68_3 & bh793_w68_4 & bh793_w68_5;
   Compressor_6_3_F200_uid1088_uid1155: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1155_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1155_Out0_copy1156);
   Compressor_6_3_F200_uid1088_bh793_uid1155_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1155_Out0_copy1156; -- output copy to hold a pipeline register if needed

   bh793_w68_12 <= Compressor_6_3_F200_uid1088_bh793_uid1155_Out0(0);
   bh793_w69_9 <= Compressor_6_3_F200_uid1088_bh793_uid1155_Out0(1);
   bh793_w70_8 <= Compressor_6_3_F200_uid1088_bh793_uid1155_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1157_In0 <= "" & bh793_w68_6 & bh793_w68_7 & bh793_w68_8;
   Compressor_23_3_F200_uid1032_bh793_uid1157_In1 <= "" & bh793_w69_0 & bh793_w69_1;
   Compressor_23_3_F200_uid1032_uid1157: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1157_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1157_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1157_Out0_copy1158);
   Compressor_23_3_F200_uid1032_bh793_uid1157_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1157_Out0_copy1158; -- output copy to hold a pipeline register if needed

   bh793_w68_13 <= Compressor_23_3_F200_uid1032_bh793_uid1157_Out0(0);
   bh793_w69_10 <= Compressor_23_3_F200_uid1032_bh793_uid1157_Out0(1);
   bh793_w70_9 <= Compressor_23_3_F200_uid1032_bh793_uid1157_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1159_In0 <= "" & bh793_w69_2 & bh793_w69_3 & bh793_w69_4 & bh793_w69_5 & bh793_w69_6 & bh793_w69_7;
   Compressor_6_3_F200_uid1088_uid1159: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1159_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1159_Out0_copy1160);
   Compressor_6_3_F200_uid1088_bh793_uid1159_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1159_Out0_copy1160; -- output copy to hold a pipeline register if needed

   bh793_w69_11 <= Compressor_6_3_F200_uid1088_bh793_uid1159_Out0(0);
   bh793_w70_10 <= Compressor_6_3_F200_uid1088_bh793_uid1159_Out0(1);
   bh793_w71_9 <= Compressor_6_3_F200_uid1088_bh793_uid1159_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1161_In0 <= "" & bh793_w70_0 & bh793_w70_1 & bh793_w70_2 & bh793_w70_3 & bh793_w70_4 & "0";
   Compressor_6_3_F200_uid1088_uid1161: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1161_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1161_Out0_copy1162);
   Compressor_6_3_F200_uid1088_bh793_uid1161_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1161_Out0_copy1162; -- output copy to hold a pipeline register if needed

   bh793_w70_11 <= Compressor_6_3_F200_uid1088_bh793_uid1161_Out0(0);
   bh793_w71_10 <= Compressor_6_3_F200_uid1088_bh793_uid1161_Out0(1);
   bh793_w72_8 <= Compressor_6_3_F200_uid1088_bh793_uid1161_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1163_In0 <= "" & bh793_w70_5 & bh793_w70_6 & bh793_w70_7;
   Compressor_3_2_F200_uid1040_uid1163: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1163_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1163_Out0_copy1164);
   Compressor_3_2_F200_uid1040_bh793_uid1163_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1163_Out0_copy1164; -- output copy to hold a pipeline register if needed

   bh793_w70_12 <= Compressor_3_2_F200_uid1040_bh793_uid1163_Out0(0);
   bh793_w71_11 <= Compressor_3_2_F200_uid1040_bh793_uid1163_Out0(1);

   Compressor_6_3_F200_uid1088_bh793_uid1165_In0 <= "" & bh793_w71_0 & bh793_w71_1 & bh793_w71_2 & bh793_w71_3 & bh793_w71_4 & bh793_w71_5;
   Compressor_6_3_F200_uid1088_uid1165: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1165_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1165_Out0_copy1166);
   Compressor_6_3_F200_uid1088_bh793_uid1165_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1165_Out0_copy1166; -- output copy to hold a pipeline register if needed

   bh793_w71_12 <= Compressor_6_3_F200_uid1088_bh793_uid1165_Out0(0);
   bh793_w72_9 <= Compressor_6_3_F200_uid1088_bh793_uid1165_Out0(1);
   bh793_w73_8 <= Compressor_6_3_F200_uid1088_bh793_uid1165_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1167_In0 <= "" & bh793_w71_6 & bh793_w71_7 & bh793_w71_8;
   Compressor_23_3_F200_uid1032_bh793_uid1167_In1 <= "" & bh793_w72_0 & bh793_w72_1;
   Compressor_23_3_F200_uid1032_uid1167: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1167_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1167_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1167_Out0_copy1168);
   Compressor_23_3_F200_uid1032_bh793_uid1167_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1167_Out0_copy1168; -- output copy to hold a pipeline register if needed

   bh793_w71_13 <= Compressor_23_3_F200_uid1032_bh793_uid1167_Out0(0);
   bh793_w72_10 <= Compressor_23_3_F200_uid1032_bh793_uid1167_Out0(1);
   bh793_w73_9 <= Compressor_23_3_F200_uid1032_bh793_uid1167_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1169_In0 <= "" & bh793_w72_2 & bh793_w72_3 & bh793_w72_4 & bh793_w72_5 & bh793_w72_6 & bh793_w72_7;
   Compressor_6_3_F200_uid1088_uid1169: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1169_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1169_Out0_copy1170);
   Compressor_6_3_F200_uid1088_bh793_uid1169_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1169_Out0_copy1170; -- output copy to hold a pipeline register if needed

   bh793_w72_11 <= Compressor_6_3_F200_uid1088_bh793_uid1169_Out0(0);
   bh793_w73_10 <= Compressor_6_3_F200_uid1088_bh793_uid1169_Out0(1);
   bh793_w74_9 <= Compressor_6_3_F200_uid1088_bh793_uid1169_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1171_In0 <= "" & bh793_w73_0 & bh793_w73_1 & bh793_w73_2 & bh793_w73_3 & bh793_w73_4 & "0";
   Compressor_6_3_F200_uid1088_uid1171: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1171_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1171_Out0_copy1172);
   Compressor_6_3_F200_uid1088_bh793_uid1171_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1171_Out0_copy1172; -- output copy to hold a pipeline register if needed

   bh793_w73_11 <= Compressor_6_3_F200_uid1088_bh793_uid1171_Out0(0);
   bh793_w74_10 <= Compressor_6_3_F200_uid1088_bh793_uid1171_Out0(1);
   bh793_w75_8 <= Compressor_6_3_F200_uid1088_bh793_uid1171_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1173_In0 <= "" & bh793_w73_5 & bh793_w73_6 & bh793_w73_7;
   Compressor_3_2_F200_uid1040_uid1173: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1173_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1173_Out0_copy1174);
   Compressor_3_2_F200_uid1040_bh793_uid1173_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1173_Out0_copy1174; -- output copy to hold a pipeline register if needed

   bh793_w73_12 <= Compressor_3_2_F200_uid1040_bh793_uid1173_Out0(0);
   bh793_w74_11 <= Compressor_3_2_F200_uid1040_bh793_uid1173_Out0(1);

   Compressor_6_3_F200_uid1088_bh793_uid1175_In0 <= "" & bh793_w74_0 & bh793_w74_1 & bh793_w74_2 & bh793_w74_3 & bh793_w74_4 & bh793_w74_5;
   Compressor_6_3_F200_uid1088_uid1175: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1175_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1175_Out0_copy1176);
   Compressor_6_3_F200_uid1088_bh793_uid1175_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1175_Out0_copy1176; -- output copy to hold a pipeline register if needed

   bh793_w74_12 <= Compressor_6_3_F200_uid1088_bh793_uid1175_Out0(0);
   bh793_w75_9 <= Compressor_6_3_F200_uid1088_bh793_uid1175_Out0(1);
   bh793_w76_8 <= Compressor_6_3_F200_uid1088_bh793_uid1175_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1177_In0 <= "" & bh793_w74_6 & bh793_w74_7 & bh793_w74_8;
   Compressor_23_3_F200_uid1032_bh793_uid1177_In1 <= "" & bh793_w75_0 & bh793_w75_1;
   Compressor_23_3_F200_uid1032_uid1177: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1177_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1177_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1177_Out0_copy1178);
   Compressor_23_3_F200_uid1032_bh793_uid1177_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1177_Out0_copy1178; -- output copy to hold a pipeline register if needed

   bh793_w74_13 <= Compressor_23_3_F200_uid1032_bh793_uid1177_Out0(0);
   bh793_w75_10 <= Compressor_23_3_F200_uid1032_bh793_uid1177_Out0(1);
   bh793_w76_9 <= Compressor_23_3_F200_uid1032_bh793_uid1177_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1179_In0 <= "" & bh793_w75_2 & bh793_w75_3 & bh793_w75_4 & bh793_w75_5 & bh793_w75_6 & bh793_w75_7;
   Compressor_6_3_F200_uid1088_uid1179: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1179_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1179_Out0_copy1180);
   Compressor_6_3_F200_uid1088_bh793_uid1179_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1179_Out0_copy1180; -- output copy to hold a pipeline register if needed

   bh793_w75_11 <= Compressor_6_3_F200_uid1088_bh793_uid1179_Out0(0);
   bh793_w76_10 <= Compressor_6_3_F200_uid1088_bh793_uid1179_Out0(1);
   bh793_w77_8 <= Compressor_6_3_F200_uid1088_bh793_uid1179_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1181_In0 <= "" & bh793_w76_0 & bh793_w76_1 & bh793_w76_2 & bh793_w76_3 & bh793_w76_4 & "0";
   Compressor_6_3_F200_uid1088_uid1181: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1181_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1181_Out0_copy1182);
   Compressor_6_3_F200_uid1088_bh793_uid1181_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1181_Out0_copy1182; -- output copy to hold a pipeline register if needed

   bh793_w76_11 <= Compressor_6_3_F200_uid1088_bh793_uid1181_Out0(0);
   bh793_w77_9 <= Compressor_6_3_F200_uid1088_bh793_uid1181_Out0(1);
   bh793_w78_7 <= Compressor_6_3_F200_uid1088_bh793_uid1181_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1183_In0 <= "" & bh793_w76_5 & bh793_w76_6 & bh793_w76_7;
   Compressor_23_3_F200_uid1032_bh793_uid1183_In1 <= "" & bh793_w77_0 & bh793_w77_1;
   Compressor_23_3_F200_uid1032_uid1183: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1183_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1183_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1183_Out0_copy1184);
   Compressor_23_3_F200_uid1032_bh793_uid1183_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1183_Out0_copy1184; -- output copy to hold a pipeline register if needed

   bh793_w76_12 <= Compressor_23_3_F200_uid1032_bh793_uid1183_Out0(0);
   bh793_w77_10 <= Compressor_23_3_F200_uid1032_bh793_uid1183_Out0(1);
   bh793_w78_8 <= Compressor_23_3_F200_uid1032_bh793_uid1183_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1185_In0 <= "" & bh793_w77_2 & bh793_w77_3 & bh793_w77_4 & bh793_w77_5 & bh793_w77_6 & bh793_w77_7;
   Compressor_6_3_F200_uid1088_uid1185: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1185_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1185_Out0_copy1186);
   Compressor_6_3_F200_uid1088_bh793_uid1185_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1185_Out0_copy1186; -- output copy to hold a pipeline register if needed

   bh793_w77_11 <= Compressor_6_3_F200_uid1088_bh793_uid1185_Out0(0);
   bh793_w78_9 <= Compressor_6_3_F200_uid1088_bh793_uid1185_Out0(1);
   bh793_w79_7 <= Compressor_6_3_F200_uid1088_bh793_uid1185_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1187_In0 <= "" & bh793_w78_0 & bh793_w78_1 & bh793_w78_2 & bh793_w78_3 & bh793_w78_4 & bh793_w78_5;
   Compressor_6_3_F200_uid1088_uid1187: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1187_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1187_Out0_copy1188);
   Compressor_6_3_F200_uid1088_bh793_uid1187_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1187_Out0_copy1188; -- output copy to hold a pipeline register if needed

   bh793_w78_10 <= Compressor_6_3_F200_uid1088_bh793_uid1187_Out0(0);
   bh793_w79_8 <= Compressor_6_3_F200_uid1088_bh793_uid1187_Out0(1);
   bh793_w80_8 <= Compressor_6_3_F200_uid1088_bh793_uid1187_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1189_In0 <= "" & bh793_w79_0 & bh793_w79_1 & bh793_w79_2 & bh793_w79_3 & bh793_w79_4 & bh793_w79_5;
   Compressor_6_3_F200_uid1088_uid1189: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1189_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1189_Out0_copy1190);
   Compressor_6_3_F200_uid1088_bh793_uid1189_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1189_Out0_copy1190; -- output copy to hold a pipeline register if needed

   bh793_w79_9 <= Compressor_6_3_F200_uid1088_bh793_uid1189_Out0(0);
   bh793_w80_9 <= Compressor_6_3_F200_uid1088_bh793_uid1189_Out0(1);
   bh793_w81_7 <= Compressor_6_3_F200_uid1088_bh793_uid1189_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1191_In0 <= "" & bh793_w80_0 & bh793_w80_1 & bh793_w80_2 & bh793_w80_3 & "0" & "0";
   Compressor_6_3_F200_uid1088_uid1191: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1191_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1191_Out0_copy1192);
   Compressor_6_3_F200_uid1088_bh793_uid1191_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1191_Out0_copy1192; -- output copy to hold a pipeline register if needed

   bh793_w80_10 <= Compressor_6_3_F200_uid1088_bh793_uid1191_Out0(0);
   bh793_w81_8 <= Compressor_6_3_F200_uid1088_bh793_uid1191_Out0(1);
   bh793_w82_7 <= Compressor_6_3_F200_uid1088_bh793_uid1191_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1193_In0 <= "" & bh793_w80_4 & bh793_w80_5 & bh793_w80_6 & bh793_w80_7;
   Compressor_14_3_F200_uid1054_bh793_uid1193_In1 <= "" & bh793_w81_0;
   Compressor_14_3_F200_uid1054_uid1193: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1193_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1193_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1193_Out0_copy1194);
   Compressor_14_3_F200_uid1054_bh793_uid1193_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1193_Out0_copy1194; -- output copy to hold a pipeline register if needed

   bh793_w80_11 <= Compressor_14_3_F200_uid1054_bh793_uid1193_Out0(0);
   bh793_w81_9 <= Compressor_14_3_F200_uid1054_bh793_uid1193_Out0(1);
   bh793_w82_8 <= Compressor_14_3_F200_uid1054_bh793_uid1193_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1195_In0 <= "" & bh793_w81_1 & bh793_w81_2 & bh793_w81_3 & bh793_w81_4 & bh793_w81_5 & bh793_w81_6;
   Compressor_6_3_F200_uid1088_uid1195: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1195_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1195_Out0_copy1196);
   Compressor_6_3_F200_uid1088_bh793_uid1195_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1195_Out0_copy1196; -- output copy to hold a pipeline register if needed

   bh793_w81_10 <= Compressor_6_3_F200_uid1088_bh793_uid1195_Out0(0);
   bh793_w82_9 <= Compressor_6_3_F200_uid1088_bh793_uid1195_Out0(1);
   bh793_w83_7 <= Compressor_6_3_F200_uid1088_bh793_uid1195_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1197_In0 <= "" & bh793_w82_0 & bh793_w82_1 & bh793_w82_2 & bh793_w82_3 & bh793_w82_4 & bh793_w82_5;
   Compressor_6_3_F200_uid1088_uid1197: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1197_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1197_Out0_copy1198);
   Compressor_6_3_F200_uid1088_bh793_uid1197_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1197_Out0_copy1198; -- output copy to hold a pipeline register if needed

   bh793_w82_10 <= Compressor_6_3_F200_uid1088_bh793_uid1197_Out0(0);
   bh793_w83_8 <= Compressor_6_3_F200_uid1088_bh793_uid1197_Out0(1);
   bh793_w84_6 <= Compressor_6_3_F200_uid1088_bh793_uid1197_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1199_In0 <= "" & bh793_w83_0 & bh793_w83_1 & bh793_w83_2 & bh793_w83_3 & bh793_w83_4 & bh793_w83_5;
   Compressor_6_3_F200_uid1088_uid1199: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1199_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1199_Out0_copy1200);
   Compressor_6_3_F200_uid1088_bh793_uid1199_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1199_Out0_copy1200; -- output copy to hold a pipeline register if needed

   bh793_w83_9 <= Compressor_6_3_F200_uid1088_bh793_uid1199_Out0(0);
   bh793_w84_7 <= Compressor_6_3_F200_uid1088_bh793_uid1199_Out0(1);
   bh793_w85_7 <= Compressor_6_3_F200_uid1088_bh793_uid1199_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1201_In0 <= "" & bh793_w84_0 & bh793_w84_1 & bh793_w84_2 & bh793_w84_3 & bh793_w84_4 & bh793_w84_5;
   Compressor_6_3_F200_uid1088_uid1201: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1201_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1201_Out0_copy1202);
   Compressor_6_3_F200_uid1088_bh793_uid1201_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1201_Out0_copy1202; -- output copy to hold a pipeline register if needed

   bh793_w84_8 <= Compressor_6_3_F200_uid1088_bh793_uid1201_Out0(0);
   bh793_w85_8 <= Compressor_6_3_F200_uid1088_bh793_uid1201_Out0(1);
   bh793_w86_6 <= Compressor_6_3_F200_uid1088_bh793_uid1201_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1203_In0 <= "" & bh793_w85_0 & bh793_w85_1 & bh793_w85_2 & bh793_w85_3 & bh793_w85_4 & bh793_w85_5;
   Compressor_6_3_F200_uid1088_uid1203: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1203_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1203_Out0_copy1204);
   Compressor_6_3_F200_uid1088_bh793_uid1203_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1203_Out0_copy1204; -- output copy to hold a pipeline register if needed

   bh793_w85_9 <= Compressor_6_3_F200_uid1088_bh793_uid1203_Out0(0);
   bh793_w86_7 <= Compressor_6_3_F200_uid1088_bh793_uid1203_Out0(1);
   bh793_w87_6 <= Compressor_6_3_F200_uid1088_bh793_uid1203_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1205_In0 <= "" & bh793_w86_0 & bh793_w86_1 & bh793_w86_2 & bh793_w86_3 & bh793_w86_4 & bh793_w86_5;
   Compressor_6_3_F200_uid1088_uid1205: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1205_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1205_Out0_copy1206);
   Compressor_6_3_F200_uid1088_bh793_uid1205_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1205_Out0_copy1206; -- output copy to hold a pipeline register if needed

   bh793_w86_8 <= Compressor_6_3_F200_uid1088_bh793_uid1205_Out0(0);
   bh793_w87_7 <= Compressor_6_3_F200_uid1088_bh793_uid1205_Out0(1);
   bh793_w88_7 <= Compressor_6_3_F200_uid1088_bh793_uid1205_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1207_In0 <= "" & bh793_w87_0 & bh793_w87_1 & bh793_w87_2 & bh793_w87_3 & bh793_w87_4 & bh793_w87_5;
   Compressor_6_3_F200_uid1088_uid1207: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1207_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1207_Out0_copy1208);
   Compressor_6_3_F200_uid1088_bh793_uid1207_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1207_Out0_copy1208; -- output copy to hold a pipeline register if needed

   bh793_w87_8 <= Compressor_6_3_F200_uid1088_bh793_uid1207_Out0(0);
   bh793_w88_8 <= Compressor_6_3_F200_uid1088_bh793_uid1207_Out0(1);
   bh793_w89_6 <= Compressor_6_3_F200_uid1088_bh793_uid1207_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1209_In0 <= "" & bh793_w88_0 & bh793_w88_1 & bh793_w88_2 & bh793_w88_3 & bh793_w88_4 & bh793_w88_5;
   Compressor_6_3_F200_uid1088_uid1209: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1209_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1209_Out0_copy1210);
   Compressor_6_3_F200_uid1088_bh793_uid1209_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1209_Out0_copy1210; -- output copy to hold a pipeline register if needed

   bh793_w88_9 <= Compressor_6_3_F200_uid1088_bh793_uid1209_Out0(0);
   bh793_w89_7 <= Compressor_6_3_F200_uid1088_bh793_uid1209_Out0(1);
   bh793_w90_6 <= Compressor_6_3_F200_uid1088_bh793_uid1209_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1211_In0 <= "" & bh793_w89_0 & bh793_w89_1 & bh793_w89_2 & bh793_w89_3 & bh793_w89_4 & bh793_w89_5;
   Compressor_6_3_F200_uid1088_uid1211: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1211_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1211_Out0_copy1212);
   Compressor_6_3_F200_uid1088_bh793_uid1211_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1211_Out0_copy1212; -- output copy to hold a pipeline register if needed

   bh793_w89_8 <= Compressor_6_3_F200_uid1088_bh793_uid1211_Out0(0);
   bh793_w90_7 <= Compressor_6_3_F200_uid1088_bh793_uid1211_Out0(1);
   bh793_w91_7 <= Compressor_6_3_F200_uid1088_bh793_uid1211_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1213_In0 <= "" & bh793_w90_0 & bh793_w90_1 & bh793_w90_2 & bh793_w90_3 & bh793_w90_4 & bh793_w90_5;
   Compressor_6_3_F200_uid1088_uid1213: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1213_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1213_Out0_copy1214);
   Compressor_6_3_F200_uid1088_bh793_uid1213_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1213_Out0_copy1214; -- output copy to hold a pipeline register if needed

   bh793_w90_8 <= Compressor_6_3_F200_uid1088_bh793_uid1213_Out0(0);
   bh793_w91_8 <= Compressor_6_3_F200_uid1088_bh793_uid1213_Out0(1);
   bh793_w92_6 <= Compressor_6_3_F200_uid1088_bh793_uid1213_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1215_In0 <= "" & bh793_w91_0 & bh793_w91_1 & bh793_w91_2 & bh793_w91_3 & bh793_w91_4 & bh793_w91_5;
   Compressor_6_3_F200_uid1088_uid1215: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1215_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1215_Out0_copy1216);
   Compressor_6_3_F200_uid1088_bh793_uid1215_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1215_Out0_copy1216; -- output copy to hold a pipeline register if needed

   bh793_w91_9 <= Compressor_6_3_F200_uid1088_bh793_uid1215_Out0(0);
   bh793_w92_7 <= Compressor_6_3_F200_uid1088_bh793_uid1215_Out0(1);
   bh793_w93_6 <= Compressor_6_3_F200_uid1088_bh793_uid1215_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1217_In0 <= "" & bh793_w92_0 & bh793_w92_1 & bh793_w92_2 & bh793_w92_3 & bh793_w92_4 & bh793_w92_5;
   Compressor_6_3_F200_uid1088_uid1217: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1217_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1217_Out0_copy1218);
   Compressor_6_3_F200_uid1088_bh793_uid1217_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1217_Out0_copy1218; -- output copy to hold a pipeline register if needed

   bh793_w92_8 <= Compressor_6_3_F200_uid1088_bh793_uid1217_Out0(0);
   bh793_w93_7 <= Compressor_6_3_F200_uid1088_bh793_uid1217_Out0(1);
   bh793_w94_7 <= Compressor_6_3_F200_uid1088_bh793_uid1217_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1219_In0 <= "" & bh793_w93_0 & bh793_w93_1 & bh793_w93_2 & bh793_w93_3 & bh793_w93_4 & bh793_w93_5;
   Compressor_6_3_F200_uid1088_uid1219: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1219_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1219_Out0_copy1220);
   Compressor_6_3_F200_uid1088_bh793_uid1219_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1219_Out0_copy1220; -- output copy to hold a pipeline register if needed

   bh793_w93_8 <= Compressor_6_3_F200_uid1088_bh793_uid1219_Out0(0);
   bh793_w94_8 <= Compressor_6_3_F200_uid1088_bh793_uid1219_Out0(1);
   bh793_w95_6 <= Compressor_6_3_F200_uid1088_bh793_uid1219_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1221_In0 <= "" & bh793_w94_0 & bh793_w94_1 & bh793_w94_2 & bh793_w94_3 & bh793_w94_4 & bh793_w94_5;
   Compressor_6_3_F200_uid1088_uid1221: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1221_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1221_Out0_copy1222);
   Compressor_6_3_F200_uid1088_bh793_uid1221_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1221_Out0_copy1222; -- output copy to hold a pipeline register if needed

   bh793_w94_9 <= Compressor_6_3_F200_uid1088_bh793_uid1221_Out0(0);
   bh793_w95_7 <= Compressor_6_3_F200_uid1088_bh793_uid1221_Out0(1);
   bh793_w96_6 <= Compressor_6_3_F200_uid1088_bh793_uid1221_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1223_In0 <= "" & bh793_w95_0 & bh793_w95_1 & bh793_w95_2 & bh793_w95_3 & bh793_w95_4 & bh793_w95_5;
   Compressor_6_3_F200_uid1088_uid1223: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1223_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1223_Out0_copy1224);
   Compressor_6_3_F200_uid1088_bh793_uid1223_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1223_Out0_copy1224; -- output copy to hold a pipeline register if needed

   bh793_w95_8 <= Compressor_6_3_F200_uid1088_bh793_uid1223_Out0(0);
   bh793_w96_7 <= Compressor_6_3_F200_uid1088_bh793_uid1223_Out0(1);
   bh793_w97_7 <= Compressor_6_3_F200_uid1088_bh793_uid1223_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1225_In0 <= "" & bh793_w96_0 & bh793_w96_1 & bh793_w96_2 & bh793_w96_3 & bh793_w96_4 & bh793_w96_5;
   Compressor_6_3_F200_uid1088_uid1225: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1225_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1225_Out0_copy1226);
   Compressor_6_3_F200_uid1088_bh793_uid1225_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1225_Out0_copy1226; -- output copy to hold a pipeline register if needed

   bh793_w96_8 <= Compressor_6_3_F200_uid1088_bh793_uid1225_Out0(0);
   bh793_w97_8 <= Compressor_6_3_F200_uid1088_bh793_uid1225_Out0(1);
   bh793_w98_6 <= Compressor_6_3_F200_uid1088_bh793_uid1225_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1227_In0 <= "" & bh793_w97_0 & bh793_w97_1 & bh793_w97_2 & bh793_w97_3 & bh793_w97_4 & bh793_w97_5;
   Compressor_6_3_F200_uid1088_uid1227: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1227_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1227_Out0_copy1228);
   Compressor_6_3_F200_uid1088_bh793_uid1227_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1227_Out0_copy1228; -- output copy to hold a pipeline register if needed

   bh793_w97_9 <= Compressor_6_3_F200_uid1088_bh793_uid1227_Out0(0);
   bh793_w98_7 <= Compressor_6_3_F200_uid1088_bh793_uid1227_Out0(1);
   bh793_w99_6 <= Compressor_6_3_F200_uid1088_bh793_uid1227_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1229_In0 <= "" & bh793_w98_0 & bh793_w98_1 & bh793_w98_2 & bh793_w98_3 & bh793_w98_4 & bh793_w98_5;
   Compressor_6_3_F200_uid1088_uid1229: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1229_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1229_Out0_copy1230);
   Compressor_6_3_F200_uid1088_bh793_uid1229_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1229_Out0_copy1230; -- output copy to hold a pipeline register if needed

   bh793_w98_8 <= Compressor_6_3_F200_uid1088_bh793_uid1229_Out0(0);
   bh793_w99_7 <= Compressor_6_3_F200_uid1088_bh793_uid1229_Out0(1);
   bh793_w100_6 <= Compressor_6_3_F200_uid1088_bh793_uid1229_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1231_In0 <= "" & bh793_w99_0 & bh793_w99_1 & bh793_w99_2 & bh793_w99_3 & bh793_w99_4 & bh793_w99_5;
   Compressor_6_3_F200_uid1088_uid1231: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1231_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1231_Out0_copy1232);
   Compressor_6_3_F200_uid1088_bh793_uid1231_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1231_Out0_copy1232; -- output copy to hold a pipeline register if needed

   bh793_w99_8 <= Compressor_6_3_F200_uid1088_bh793_uid1231_Out0(0);
   bh793_w100_7 <= Compressor_6_3_F200_uid1088_bh793_uid1231_Out0(1);
   bh793_w101_3 <= Compressor_6_3_F200_uid1088_bh793_uid1231_Out0(2);

   Compressor_6_3_F200_uid1088_bh793_uid1233_In0 <= "" & bh793_w100_0 & bh793_w100_1 & bh793_w100_2 & bh793_w100_3 & bh793_w100_4 & bh793_w100_5;
   Compressor_6_3_F200_uid1088_uid1233: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1233_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1233_Out0_copy1234);
   Compressor_6_3_F200_uid1088_bh793_uid1233_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1233_Out0_copy1234; -- output copy to hold a pipeline register if needed

   bh793_w100_8 <= Compressor_6_3_F200_uid1088_bh793_uid1233_Out0(0);
   bh793_w101_4 <= Compressor_6_3_F200_uid1088_bh793_uid1233_Out0(1);
   bh793_w102_4 <= Compressor_6_3_F200_uid1088_bh793_uid1233_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1235_In0 <= "" & bh793_w101_0 & bh793_w101_1 & bh793_w101_2;
   Compressor_3_2_F200_uid1040_uid1235: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1235_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1235_Out0_copy1236);
   Compressor_3_2_F200_uid1040_bh793_uid1235_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1235_Out0_copy1236; -- output copy to hold a pipeline register if needed

   bh793_w101_5 <= Compressor_3_2_F200_uid1040_bh793_uid1235_Out0(0);
   bh793_w102_5 <= Compressor_3_2_F200_uid1040_bh793_uid1235_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1237_In0 <= "" & bh793_w102_0 & bh793_w102_1 & bh793_w102_2 & bh793_w102_3;
   Compressor_14_3_F200_uid1054_bh793_uid1237_In1 <= "" & bh793_w103_0;
   Compressor_14_3_F200_uid1054_uid1237: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1237_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1237_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1237_Out0_copy1238);
   Compressor_14_3_F200_uid1054_bh793_uid1237_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1237_Out0_copy1238; -- output copy to hold a pipeline register if needed

   bh793_w102_6 <= Compressor_14_3_F200_uid1054_bh793_uid1237_Out0(0);
   bh793_w103_2 <= Compressor_14_3_F200_uid1054_bh793_uid1237_Out0(1);
   bh793_w104_1 <= Compressor_14_3_F200_uid1054_bh793_uid1237_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1239_In0 <= "" & bh793_w19_3 & bh793_w19_2 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1239_In1 <= "" & bh793_w20_2;
   Compressor_14_3_F200_uid1054_uid1239: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1239_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1239_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1239_Out0_copy1240);
   Compressor_14_3_F200_uid1054_bh793_uid1239_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1239_Out0_copy1240; -- output copy to hold a pipeline register if needed

   bh793_w19_4 <= Compressor_14_3_F200_uid1054_bh793_uid1239_Out0(0);
   bh793_w20_3 <= Compressor_14_3_F200_uid1054_bh793_uid1239_Out0(1);
   bh793_w21_4 <= Compressor_14_3_F200_uid1054_bh793_uid1239_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1241_In0 <= "" & bh793_w21_3 & bh793_w21_2 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1241_In1 <= "" & bh793_w22_2;
   Compressor_14_3_F200_uid1054_uid1241: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1241_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1241_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1241_Out0_copy1242);
   Compressor_14_3_F200_uid1054_bh793_uid1241_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1241_Out0_copy1242; -- output copy to hold a pipeline register if needed

   bh793_w21_5 <= Compressor_14_3_F200_uid1054_bh793_uid1241_Out0(0);
   bh793_w22_3 <= Compressor_14_3_F200_uid1054_bh793_uid1241_Out0(1);
   bh793_w23_4 <= Compressor_14_3_F200_uid1054_bh793_uid1241_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1243_In0 <= "" & bh793_w23_3 & bh793_w23_2 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1243_In1 <= "" & bh793_w24_4 & bh793_w24_3;
   Compressor_23_3_F200_uid1032_uid1243: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1243_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1243_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1243_Out0_copy1244);
   Compressor_23_3_F200_uid1032_bh793_uid1243_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1243_Out0_copy1244; -- output copy to hold a pipeline register if needed

   bh793_w23_5 <= Compressor_23_3_F200_uid1032_bh793_uid1243_Out0(0);
   bh793_w24_5 <= Compressor_23_3_F200_uid1032_bh793_uid1243_Out0(1);
   bh793_w25_4 <= Compressor_23_3_F200_uid1032_bh793_uid1243_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1245_In0 <= "" & bh793_w25_2 & bh793_w25_3 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1245_In1 <= "" & bh793_w26_4 & bh793_w26_3;
   Compressor_23_3_F200_uid1032_uid1245: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1245_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1245_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1245_Out0_copy1246);
   Compressor_23_3_F200_uid1032_bh793_uid1245_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1245_Out0_copy1246; -- output copy to hold a pipeline register if needed

   bh793_w25_5 <= Compressor_23_3_F200_uid1032_bh793_uid1245_Out0(0);
   bh793_w26_5 <= Compressor_23_3_F200_uid1032_bh793_uid1245_Out0(1);
   bh793_w27_4 <= Compressor_23_3_F200_uid1032_bh793_uid1245_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1247_In0 <= "" & bh793_w27_2 & bh793_w27_3 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1247_In1 <= "" & bh793_w28_4 & bh793_w28_3;
   Compressor_23_3_F200_uid1032_uid1247: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1247_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1247_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1247_Out0_copy1248);
   Compressor_23_3_F200_uid1032_bh793_uid1247_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1247_Out0_copy1248; -- output copy to hold a pipeline register if needed

   bh793_w27_5 <= Compressor_23_3_F200_uid1032_bh793_uid1247_Out0(0);
   bh793_w28_5 <= Compressor_23_3_F200_uid1032_bh793_uid1247_Out0(1);
   bh793_w29_4 <= Compressor_23_3_F200_uid1032_bh793_uid1247_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1249_In0 <= "" & bh793_w29_2 & bh793_w29_3 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1249_In1 <= "" & bh793_w30_4 & bh793_w30_3;
   Compressor_23_3_F200_uid1032_uid1249: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1249_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1249_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1249_Out0_copy1250);
   Compressor_23_3_F200_uid1032_bh793_uid1249_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1249_Out0_copy1250; -- output copy to hold a pipeline register if needed

   bh793_w29_5 <= Compressor_23_3_F200_uid1032_bh793_uid1249_Out0(0);
   bh793_w30_5 <= Compressor_23_3_F200_uid1032_bh793_uid1249_Out0(1);
   bh793_w31_4 <= Compressor_23_3_F200_uid1032_bh793_uid1249_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1251_In0 <= "" & bh793_w31_2 & bh793_w31_3 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1251_In1 <= "" & bh793_w32_4 & bh793_w32_3;
   Compressor_23_3_F200_uid1032_uid1251: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1251_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1251_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1251_Out0_copy1252);
   Compressor_23_3_F200_uid1032_bh793_uid1251_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1251_Out0_copy1252; -- output copy to hold a pipeline register if needed

   bh793_w31_5 <= Compressor_23_3_F200_uid1032_bh793_uid1251_Out0(0);
   bh793_w32_5 <= Compressor_23_3_F200_uid1032_bh793_uid1251_Out0(1);
   bh793_w33_4 <= Compressor_23_3_F200_uid1032_bh793_uid1251_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1253_In0 <= "" & bh793_w33_2 & bh793_w33_3 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1253_In1 <= "" & bh793_w34_5 & bh793_w34_4;
   Compressor_23_3_F200_uid1032_uid1253: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1253_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1253_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1253_Out0_copy1254);
   Compressor_23_3_F200_uid1032_bh793_uid1253_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1253_Out0_copy1254; -- output copy to hold a pipeline register if needed

   bh793_w33_5 <= Compressor_23_3_F200_uid1032_bh793_uid1253_Out0(0);
   bh793_w34_6 <= Compressor_23_3_F200_uid1032_bh793_uid1253_Out0(1);
   bh793_w35_6 <= Compressor_23_3_F200_uid1032_bh793_uid1253_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1255_In0 <= "" & bh793_w35_5 & bh793_w35_4 & "0";
   Compressor_3_2_F200_uid1040_uid1255: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1255_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1255_Out0_copy1256);
   Compressor_3_2_F200_uid1040_bh793_uid1255_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1255_Out0_copy1256; -- output copy to hold a pipeline register if needed

   bh793_w35_7 <= Compressor_3_2_F200_uid1040_bh793_uid1255_Out0(0);
   bh793_w36_7 <= Compressor_3_2_F200_uid1040_bh793_uid1255_Out0(1);

   Compressor_23_3_F200_uid1032_bh793_uid1257_In0 <= "" & bh793_w36_6 & bh793_w36_5 & bh793_w36_4;
   Compressor_23_3_F200_uid1032_bh793_uid1257_In1 <= "" & bh793_w37_5 & bh793_w37_4;
   Compressor_23_3_F200_uid1032_uid1257: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1257_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1257_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1257_Out0_copy1258);
   Compressor_23_3_F200_uid1032_bh793_uid1257_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1257_Out0_copy1258; -- output copy to hold a pipeline register if needed

   bh793_w36_8 <= Compressor_23_3_F200_uid1032_bh793_uid1257_Out0(0);
   bh793_w37_6 <= Compressor_23_3_F200_uid1032_bh793_uid1257_Out0(1);
   bh793_w38_7 <= Compressor_23_3_F200_uid1032_bh793_uid1257_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1259_In0 <= "" & bh793_w38_6 & bh793_w38_5 & bh793_w38_4;
   Compressor_23_3_F200_uid1032_bh793_uid1259_In1 <= "" & bh793_w39_5 & bh793_w39_4;
   Compressor_23_3_F200_uid1032_uid1259: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1259_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1259_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1259_Out0_copy1260);
   Compressor_23_3_F200_uid1032_bh793_uid1259_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1259_Out0_copy1260; -- output copy to hold a pipeline register if needed

   bh793_w38_8 <= Compressor_23_3_F200_uid1032_bh793_uid1259_Out0(0);
   bh793_w39_6 <= Compressor_23_3_F200_uid1032_bh793_uid1259_Out0(1);
   bh793_w40_7 <= Compressor_23_3_F200_uid1032_bh793_uid1259_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1261_In0 <= "" & bh793_w40_6 & bh793_w40_5 & bh793_w40_4;
   Compressor_23_3_F200_uid1032_bh793_uid1261_In1 <= "" & bh793_w41_5 & bh793_w41_4;
   Compressor_23_3_F200_uid1032_uid1261: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1261_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1261_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1261_Out0_copy1262);
   Compressor_23_3_F200_uid1032_bh793_uid1261_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1261_Out0_copy1262; -- output copy to hold a pipeline register if needed

   bh793_w40_8 <= Compressor_23_3_F200_uid1032_bh793_uid1261_Out0(0);
   bh793_w41_6 <= Compressor_23_3_F200_uid1032_bh793_uid1261_Out0(1);
   bh793_w42_7 <= Compressor_23_3_F200_uid1032_bh793_uid1261_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1263_In0 <= "" & bh793_w42_6 & bh793_w42_5 & bh793_w42_4;
   Compressor_23_3_F200_uid1032_bh793_uid1263_In1 <= "" & bh793_w43_5 & bh793_w43_4;
   Compressor_23_3_F200_uid1032_uid1263: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1263_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1263_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1263_Out0_copy1264);
   Compressor_23_3_F200_uid1032_bh793_uid1263_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1263_Out0_copy1264; -- output copy to hold a pipeline register if needed

   bh793_w42_8 <= Compressor_23_3_F200_uid1032_bh793_uid1263_Out0(0);
   bh793_w43_6 <= Compressor_23_3_F200_uid1032_bh793_uid1263_Out0(1);
   bh793_w44_7 <= Compressor_23_3_F200_uid1032_bh793_uid1263_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1265_In0 <= "" & bh793_w44_6 & bh793_w44_5 & bh793_w44_4;
   Compressor_23_3_F200_uid1032_bh793_uid1265_In1 <= "" & bh793_w45_5 & bh793_w45_4;
   Compressor_23_3_F200_uid1032_uid1265: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1265_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1265_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1265_Out0_copy1266);
   Compressor_23_3_F200_uid1032_bh793_uid1265_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1265_Out0_copy1266; -- output copy to hold a pipeline register if needed

   bh793_w44_8 <= Compressor_23_3_F200_uid1032_bh793_uid1265_Out0(0);
   bh793_w45_6 <= Compressor_23_3_F200_uid1032_bh793_uid1265_Out0(1);
   bh793_w46_7 <= Compressor_23_3_F200_uid1032_bh793_uid1265_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1267_In0 <= "" & bh793_w46_6 & bh793_w46_5 & bh793_w46_4;
   Compressor_23_3_F200_uid1032_bh793_uid1267_In1 <= "" & bh793_w47_5 & bh793_w47_4;
   Compressor_23_3_F200_uid1032_uid1267: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1267_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1267_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1267_Out0_copy1268);
   Compressor_23_3_F200_uid1032_bh793_uid1267_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1267_Out0_copy1268; -- output copy to hold a pipeline register if needed

   bh793_w46_8 <= Compressor_23_3_F200_uid1032_bh793_uid1267_Out0(0);
   bh793_w47_6 <= Compressor_23_3_F200_uid1032_bh793_uid1267_Out0(1);
   bh793_w48_8 <= Compressor_23_3_F200_uid1032_bh793_uid1267_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1269_In0 <= "" & bh793_w48_7 & bh793_w48_6 & bh793_w48_5 & bh793_w48_4;
   Compressor_14_3_F200_uid1054_bh793_uid1269_In1 <= "" & "0";
   Compressor_14_3_F200_uid1054_uid1269: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1269_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1269_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1269_Out0_copy1270);
   Compressor_14_3_F200_uid1054_bh793_uid1269_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1269_Out0_copy1270; -- output copy to hold a pipeline register if needed

   bh793_w48_9 <= Compressor_14_3_F200_uid1054_bh793_uid1269_Out0(0);
   bh793_w49_7 <= Compressor_14_3_F200_uid1054_bh793_uid1269_Out0(1);
   bh793_w50_9 <= Compressor_14_3_F200_uid1054_bh793_uid1269_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1271_In0 <= "" & bh793_w49_6 & bh793_w49_5 & bh793_w49_4;
   Compressor_3_2_F200_uid1040_uid1271: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1271_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1271_Out0_copy1272);
   Compressor_3_2_F200_uid1040_bh793_uid1271_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1271_Out0_copy1272; -- output copy to hold a pipeline register if needed

   bh793_w49_8 <= Compressor_3_2_F200_uid1040_bh793_uid1271_Out0(0);
   bh793_w50_10 <= Compressor_3_2_F200_uid1040_bh793_uid1271_Out0(1);

   Compressor_23_3_F200_uid1032_bh793_uid1273_In0 <= "" & bh793_w50_8 & bh793_w50_7 & bh793_w50_6;
   Compressor_23_3_F200_uid1032_bh793_uid1273_In1 <= "" & bh793_w51_10 & bh793_w51_9;
   Compressor_23_3_F200_uid1032_uid1273: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1273_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1273_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1273_Out0_copy1274);
   Compressor_23_3_F200_uid1032_bh793_uid1273_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1273_Out0_copy1274; -- output copy to hold a pipeline register if needed

   bh793_w50_11 <= Compressor_23_3_F200_uid1032_bh793_uid1273_Out0(0);
   bh793_w51_11 <= Compressor_23_3_F200_uid1032_bh793_uid1273_Out0(1);
   bh793_w52_14 <= Compressor_23_3_F200_uid1032_bh793_uid1273_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1275_In0 <= "" & bh793_w52_13 & bh793_w52_12 & bh793_w52_11 & bh793_w52_10;
   Compressor_14_3_F200_uid1054_bh793_uid1275_In1 <= "" & bh793_w53_12;
   Compressor_14_3_F200_uid1054_uid1275: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1275_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1275_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1275_Out0_copy1276);
   Compressor_14_3_F200_uid1054_bh793_uid1275_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1275_Out0_copy1276; -- output copy to hold a pipeline register if needed

   bh793_w52_15 <= Compressor_14_3_F200_uid1054_bh793_uid1275_Out0(0);
   bh793_w53_13 <= Compressor_14_3_F200_uid1054_bh793_uid1275_Out0(1);
   bh793_w54_15 <= Compressor_14_3_F200_uid1054_bh793_uid1275_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1277_In0 <= "" & bh793_w53_11 & bh793_w53_10 & bh793_w53_9 & bh793_w53_8;
   Compressor_14_3_F200_uid1054_bh793_uid1277_In1 <= "" & bh793_w54_14;
   Compressor_14_3_F200_uid1054_uid1277: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1277_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1277_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1277_Out0_copy1278);
   Compressor_14_3_F200_uid1054_bh793_uid1277_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1277_Out0_copy1278; -- output copy to hold a pipeline register if needed

   bh793_w53_14 <= Compressor_14_3_F200_uid1054_bh793_uid1277_Out0(0);
   bh793_w54_16 <= Compressor_14_3_F200_uid1054_bh793_uid1277_Out0(1);
   bh793_w55_14 <= Compressor_14_3_F200_uid1054_bh793_uid1277_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1279_In0 <= "" & bh793_w54_13 & bh793_w54_12 & bh793_w54_11 & bh793_w54_10;
   Compressor_14_3_F200_uid1054_bh793_uid1279_In1 <= "" & bh793_w55_11;
   Compressor_14_3_F200_uid1054_uid1279: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1279_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1279_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1279_Out0_copy1280);
   Compressor_14_3_F200_uid1054_bh793_uid1279_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1279_Out0_copy1280; -- output copy to hold a pipeline register if needed

   bh793_w54_17 <= Compressor_14_3_F200_uid1054_bh793_uid1279_Out0(0);
   bh793_w55_15 <= Compressor_14_3_F200_uid1054_bh793_uid1279_Out0(1);
   bh793_w56_15 <= Compressor_14_3_F200_uid1054_bh793_uid1279_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1281_In0 <= "" & bh793_w55_13 & bh793_w55_12 & bh793_w55_10;
   Compressor_3_2_F200_uid1040_uid1281: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1281_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1281_Out0_copy1282);
   Compressor_3_2_F200_uid1040_bh793_uid1281_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1281_Out0_copy1282; -- output copy to hold a pipeline register if needed

   bh793_w55_16 <= Compressor_3_2_F200_uid1040_bh793_uid1281_Out0(0);
   bh793_w56_16 <= Compressor_3_2_F200_uid1040_bh793_uid1281_Out0(1);

   Compressor_6_3_F200_uid1088_bh793_uid1283_In0 <= "" & bh793_w56_10 & bh793_w56_14 & bh793_w56_13 & bh793_w56_12 & bh793_w56_11 & bh793_w56_9;
   Compressor_6_3_F200_uid1088_uid1283: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1283_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1283_Out0_copy1284);
   Compressor_6_3_F200_uid1088_bh793_uid1283_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1283_Out0_copy1284; -- output copy to hold a pipeline register if needed

   bh793_w56_17 <= Compressor_6_3_F200_uid1088_bh793_uid1283_Out0(0);
   bh793_w57_15 <= Compressor_6_3_F200_uid1088_bh793_uid1283_Out0(1);
   bh793_w58_14 <= Compressor_6_3_F200_uid1088_bh793_uid1283_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1285_In0 <= "" & bh793_w57_14 & bh793_w57_13 & bh793_w57_12 & bh793_w57_11;
   Compressor_14_3_F200_uid1054_bh793_uid1285_In1 <= "" & bh793_w58_11;
   Compressor_14_3_F200_uid1054_uid1285: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1285_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1285_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1285_Out0_copy1286);
   Compressor_14_3_F200_uid1054_bh793_uid1285_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1285_Out0_copy1286; -- output copy to hold a pipeline register if needed

   bh793_w57_16 <= Compressor_14_3_F200_uid1054_bh793_uid1285_Out0(0);
   bh793_w58_15 <= Compressor_14_3_F200_uid1054_bh793_uid1285_Out0(1);
   bh793_w59_15 <= Compressor_14_3_F200_uid1054_bh793_uid1285_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1287_In0 <= "" & bh793_w58_13 & bh793_w58_12 & bh793_w58_10;
   Compressor_3_2_F200_uid1040_uid1287: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1287_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1287_Out0_copy1288);
   Compressor_3_2_F200_uid1040_bh793_uid1287_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1287_Out0_copy1288; -- output copy to hold a pipeline register if needed

   bh793_w58_16 <= Compressor_3_2_F200_uid1040_bh793_uid1287_Out0(0);
   bh793_w59_16 <= Compressor_3_2_F200_uid1040_bh793_uid1287_Out0(1);

   Compressor_6_3_F200_uid1088_bh793_uid1289_In0 <= "" & bh793_w59_10 & bh793_w59_14 & bh793_w59_13 & bh793_w59_12 & bh793_w59_11 & bh793_w59_9;
   Compressor_6_3_F200_uid1088_uid1289: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1289_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1289_Out0_copy1290);
   Compressor_6_3_F200_uid1088_bh793_uid1289_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1289_Out0_copy1290; -- output copy to hold a pipeline register if needed

   bh793_w59_17 <= Compressor_6_3_F200_uid1088_bh793_uid1289_Out0(0);
   bh793_w60_15 <= Compressor_6_3_F200_uid1088_bh793_uid1289_Out0(1);
   bh793_w61_14 <= Compressor_6_3_F200_uid1088_bh793_uid1289_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1291_In0 <= "" & bh793_w60_14 & bh793_w60_13 & bh793_w60_12 & bh793_w60_11;
   Compressor_14_3_F200_uid1054_bh793_uid1291_In1 <= "" & bh793_w61_11;
   Compressor_14_3_F200_uid1054_uid1291: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1291_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1291_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1291_Out0_copy1292);
   Compressor_14_3_F200_uid1054_bh793_uid1291_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1291_Out0_copy1292; -- output copy to hold a pipeline register if needed

   bh793_w60_16 <= Compressor_14_3_F200_uid1054_bh793_uid1291_Out0(0);
   bh793_w61_15 <= Compressor_14_3_F200_uid1054_bh793_uid1291_Out0(1);
   bh793_w62_15 <= Compressor_14_3_F200_uid1054_bh793_uid1291_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1293_In0 <= "" & bh793_w61_13 & bh793_w61_12 & bh793_w61_10;
   Compressor_3_2_F200_uid1040_uid1293: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1293_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1293_Out0_copy1294);
   Compressor_3_2_F200_uid1040_bh793_uid1293_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1293_Out0_copy1294; -- output copy to hold a pipeline register if needed

   bh793_w61_16 <= Compressor_3_2_F200_uid1040_bh793_uid1293_Out0(0);
   bh793_w62_16 <= Compressor_3_2_F200_uid1040_bh793_uid1293_Out0(1);

   Compressor_6_3_F200_uid1088_bh793_uid1295_In0 <= "" & bh793_w62_10 & bh793_w62_14 & bh793_w62_13 & bh793_w62_12 & bh793_w62_11 & bh793_w62_9;
   Compressor_6_3_F200_uid1088_uid1295: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1295_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1295_Out0_copy1296);
   Compressor_6_3_F200_uid1088_bh793_uid1295_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1295_Out0_copy1296; -- output copy to hold a pipeline register if needed

   bh793_w62_17 <= Compressor_6_3_F200_uid1088_bh793_uid1295_Out0(0);
   bh793_w63_15 <= Compressor_6_3_F200_uid1088_bh793_uid1295_Out0(1);
   bh793_w64_14 <= Compressor_6_3_F200_uid1088_bh793_uid1295_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1297_In0 <= "" & bh793_w63_14 & bh793_w63_13 & bh793_w63_12 & bh793_w63_11;
   Compressor_14_3_F200_uid1054_bh793_uid1297_In1 <= "" & bh793_w64_11;
   Compressor_14_3_F200_uid1054_uid1297: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1297_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1297_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1297_Out0_copy1298);
   Compressor_14_3_F200_uid1054_bh793_uid1297_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1297_Out0_copy1298; -- output copy to hold a pipeline register if needed

   bh793_w63_16 <= Compressor_14_3_F200_uid1054_bh793_uid1297_Out0(0);
   bh793_w64_15 <= Compressor_14_3_F200_uid1054_bh793_uid1297_Out0(1);
   bh793_w65_15 <= Compressor_14_3_F200_uid1054_bh793_uid1297_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1299_In0 <= "" & bh793_w64_13 & bh793_w64_12 & bh793_w64_10;
   Compressor_3_2_F200_uid1040_uid1299: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1299_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1299_Out0_copy1300);
   Compressor_3_2_F200_uid1040_bh793_uid1299_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1299_Out0_copy1300; -- output copy to hold a pipeline register if needed

   bh793_w64_16 <= Compressor_3_2_F200_uid1040_bh793_uid1299_Out0(0);
   bh793_w65_16 <= Compressor_3_2_F200_uid1040_bh793_uid1299_Out0(1);

   Compressor_6_3_F200_uid1088_bh793_uid1301_In0 <= "" & bh793_w65_10 & bh793_w65_14 & bh793_w65_13 & bh793_w65_12 & bh793_w65_11 & bh793_w65_9;
   Compressor_6_3_F200_uid1088_uid1301: Compressor_6_3_F200_uid1088
      port map ( X0 => Compressor_6_3_F200_uid1088_bh793_uid1301_In0,
                 R => Compressor_6_3_F200_uid1088_bh793_uid1301_Out0_copy1302);
   Compressor_6_3_F200_uid1088_bh793_uid1301_Out0 <= Compressor_6_3_F200_uid1088_bh793_uid1301_Out0_copy1302; -- output copy to hold a pipeline register if needed

   bh793_w65_17 <= Compressor_6_3_F200_uid1088_bh793_uid1301_Out0(0);
   bh793_w66_14 <= Compressor_6_3_F200_uid1088_bh793_uid1301_Out0(1);
   bh793_w67_13 <= Compressor_6_3_F200_uid1088_bh793_uid1301_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1303_In0 <= "" & bh793_w66_11 & bh793_w66_13 & bh793_w66_12 & bh793_w66_10;
   Compressor_14_3_F200_uid1054_bh793_uid1303_In1 <= "" & bh793_w67_9;
   Compressor_14_3_F200_uid1054_uid1303: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1303_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1303_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1303_Out0_copy1304);
   Compressor_14_3_F200_uid1054_bh793_uid1303_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1303_Out0_copy1304; -- output copy to hold a pipeline register if needed

   bh793_w66_15 <= Compressor_14_3_F200_uid1054_bh793_uid1303_Out0(0);
   bh793_w67_14 <= Compressor_14_3_F200_uid1054_bh793_uid1303_Out0(1);
   bh793_w68_14 <= Compressor_14_3_F200_uid1054_bh793_uid1303_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1305_In0 <= "" & bh793_w67_12 & bh793_w67_11 & bh793_w67_10 & bh793_w67_8;
   Compressor_14_3_F200_uid1054_bh793_uid1305_In1 <= "" & bh793_w68_13;
   Compressor_14_3_F200_uid1054_uid1305: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1305_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1305_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1305_Out0_copy1306);
   Compressor_14_3_F200_uid1054_bh793_uid1305_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1305_Out0_copy1306; -- output copy to hold a pipeline register if needed

   bh793_w67_15 <= Compressor_14_3_F200_uid1054_bh793_uid1305_Out0(0);
   bh793_w68_15 <= Compressor_14_3_F200_uid1054_bh793_uid1305_Out0(1);
   bh793_w69_12 <= Compressor_14_3_F200_uid1054_bh793_uid1305_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1307_In0 <= "" & bh793_w68_12 & bh793_w68_11 & bh793_w68_10 & bh793_w68_9;
   Compressor_14_3_F200_uid1054_bh793_uid1307_In1 <= "" & bh793_w69_11;
   Compressor_14_3_F200_uid1054_uid1307: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1307_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1307_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1307_Out0_copy1308);
   Compressor_14_3_F200_uid1054_bh793_uid1307_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1307_Out0_copy1308; -- output copy to hold a pipeline register if needed

   bh793_w68_16 <= Compressor_14_3_F200_uid1054_bh793_uid1307_Out0(0);
   bh793_w69_13 <= Compressor_14_3_F200_uid1054_bh793_uid1307_Out0(1);
   bh793_w70_13 <= Compressor_14_3_F200_uid1054_bh793_uid1307_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1309_In0 <= "" & bh793_w69_10 & bh793_w69_9 & bh793_w69_8;
   Compressor_3_2_F200_uid1040_uid1309: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1309_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1309_Out0_copy1310);
   Compressor_3_2_F200_uid1040_bh793_uid1309_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1309_Out0_copy1310; -- output copy to hold a pipeline register if needed

   bh793_w69_14 <= Compressor_3_2_F200_uid1040_bh793_uid1309_Out0(0);
   bh793_w70_14 <= Compressor_3_2_F200_uid1040_bh793_uid1309_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1311_In0 <= "" & bh793_w70_12 & bh793_w70_11 & bh793_w70_10 & bh793_w70_9;
   Compressor_14_3_F200_uid1054_bh793_uid1311_In1 <= "" & bh793_w71_13;
   Compressor_14_3_F200_uid1054_uid1311: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1311_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1311_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1311_Out0_copy1312);
   Compressor_14_3_F200_uid1054_bh793_uid1311_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1311_Out0_copy1312; -- output copy to hold a pipeline register if needed

   bh793_w70_15 <= Compressor_14_3_F200_uid1054_bh793_uid1311_Out0(0);
   bh793_w71_14 <= Compressor_14_3_F200_uid1054_bh793_uid1311_Out0(1);
   bh793_w72_12 <= Compressor_14_3_F200_uid1054_bh793_uid1311_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1313_In0 <= "" & bh793_w71_12 & bh793_w71_11 & bh793_w71_10 & bh793_w71_9;
   Compressor_14_3_F200_uid1054_bh793_uid1313_In1 <= "" & bh793_w72_11;
   Compressor_14_3_F200_uid1054_uid1313: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1313_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1313_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1313_Out0_copy1314);
   Compressor_14_3_F200_uid1054_bh793_uid1313_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1313_Out0_copy1314; -- output copy to hold a pipeline register if needed

   bh793_w71_15 <= Compressor_14_3_F200_uid1054_bh793_uid1313_Out0(0);
   bh793_w72_13 <= Compressor_14_3_F200_uid1054_bh793_uid1313_Out0(1);
   bh793_w73_13 <= Compressor_14_3_F200_uid1054_bh793_uid1313_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1315_In0 <= "" & bh793_w72_10 & bh793_w72_9 & bh793_w72_8;
   Compressor_3_2_F200_uid1040_uid1315: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1315_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1315_Out0_copy1316);
   Compressor_3_2_F200_uid1040_bh793_uid1315_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1315_Out0_copy1316; -- output copy to hold a pipeline register if needed

   bh793_w72_14 <= Compressor_3_2_F200_uid1040_bh793_uid1315_Out0(0);
   bh793_w73_14 <= Compressor_3_2_F200_uid1040_bh793_uid1315_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1317_In0 <= "" & bh793_w73_12 & bh793_w73_11 & bh793_w73_10 & bh793_w73_9;
   Compressor_14_3_F200_uid1054_bh793_uid1317_In1 <= "" & bh793_w74_13;
   Compressor_14_3_F200_uid1054_uid1317: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1317_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1317_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1317_Out0_copy1318);
   Compressor_14_3_F200_uid1054_bh793_uid1317_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1317_Out0_copy1318; -- output copy to hold a pipeline register if needed

   bh793_w73_15 <= Compressor_14_3_F200_uid1054_bh793_uid1317_Out0(0);
   bh793_w74_14 <= Compressor_14_3_F200_uid1054_bh793_uid1317_Out0(1);
   bh793_w75_12 <= Compressor_14_3_F200_uid1054_bh793_uid1317_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1319_In0 <= "" & bh793_w74_12 & bh793_w74_11 & bh793_w74_10 & bh793_w74_9;
   Compressor_14_3_F200_uid1054_bh793_uid1319_In1 <= "" & bh793_w75_11;
   Compressor_14_3_F200_uid1054_uid1319: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1319_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1319_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1319_Out0_copy1320);
   Compressor_14_3_F200_uid1054_bh793_uid1319_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1319_Out0_copy1320; -- output copy to hold a pipeline register if needed

   bh793_w74_15 <= Compressor_14_3_F200_uid1054_bh793_uid1319_Out0(0);
   bh793_w75_13 <= Compressor_14_3_F200_uid1054_bh793_uid1319_Out0(1);
   bh793_w76_13 <= Compressor_14_3_F200_uid1054_bh793_uid1319_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1321_In0 <= "" & bh793_w75_10 & bh793_w75_9 & bh793_w75_8;
   Compressor_3_2_F200_uid1040_uid1321: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1321_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1321_Out0_copy1322);
   Compressor_3_2_F200_uid1040_bh793_uid1321_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1321_Out0_copy1322; -- output copy to hold a pipeline register if needed

   bh793_w75_14 <= Compressor_3_2_F200_uid1040_bh793_uid1321_Out0(0);
   bh793_w76_14 <= Compressor_3_2_F200_uid1040_bh793_uid1321_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1323_In0 <= "" & bh793_w76_12 & bh793_w76_11 & bh793_w76_10 & bh793_w76_9;
   Compressor_14_3_F200_uid1054_bh793_uid1323_In1 <= "" & bh793_w77_11;
   Compressor_14_3_F200_uid1054_uid1323: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1323_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1323_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1323_Out0_copy1324);
   Compressor_14_3_F200_uid1054_bh793_uid1323_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1323_Out0_copy1324; -- output copy to hold a pipeline register if needed

   bh793_w76_15 <= Compressor_14_3_F200_uid1054_bh793_uid1323_Out0(0);
   bh793_w77_12 <= Compressor_14_3_F200_uid1054_bh793_uid1323_Out0(1);
   bh793_w78_11 <= Compressor_14_3_F200_uid1054_bh793_uid1323_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1325_In0 <= "" & bh793_w77_10 & bh793_w77_9 & bh793_w77_8;
   Compressor_3_2_F200_uid1040_uid1325: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1325_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1325_Out0_copy1326);
   Compressor_3_2_F200_uid1040_bh793_uid1325_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1325_Out0_copy1326; -- output copy to hold a pipeline register if needed

   bh793_w77_13 <= Compressor_3_2_F200_uid1040_bh793_uid1325_Out0(0);
   bh793_w78_12 <= Compressor_3_2_F200_uid1040_bh793_uid1325_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1327_In0 <= "" & bh793_w78_10 & bh793_w78_9 & bh793_w78_8 & bh793_w78_7;
   Compressor_14_3_F200_uid1054_bh793_uid1327_In1 <= "" & bh793_w79_9;
   Compressor_14_3_F200_uid1054_uid1327: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1327_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1327_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1327_Out0_copy1328);
   Compressor_14_3_F200_uid1054_bh793_uid1327_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1327_Out0_copy1328; -- output copy to hold a pipeline register if needed

   bh793_w78_13 <= Compressor_14_3_F200_uid1054_bh793_uid1327_Out0(0);
   bh793_w79_10 <= Compressor_14_3_F200_uid1054_bh793_uid1327_Out0(1);
   bh793_w80_12 <= Compressor_14_3_F200_uid1054_bh793_uid1327_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1329_In0 <= "" & bh793_w79_8 & bh793_w79_7 & bh793_w79_6;
   Compressor_3_2_F200_uid1040_uid1329: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1329_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1329_Out0_copy1330);
   Compressor_3_2_F200_uid1040_bh793_uid1329_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1329_Out0_copy1330; -- output copy to hold a pipeline register if needed

   bh793_w79_11 <= Compressor_3_2_F200_uid1040_bh793_uid1329_Out0(0);
   bh793_w80_13 <= Compressor_3_2_F200_uid1040_bh793_uid1329_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1331_In0 <= "" & bh793_w80_11 & bh793_w80_10 & bh793_w80_9 & bh793_w80_8;
   Compressor_14_3_F200_uid1054_bh793_uid1331_In1 <= "" & bh793_w81_10;
   Compressor_14_3_F200_uid1054_uid1331: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1331_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1331_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1331_Out0_copy1332);
   Compressor_14_3_F200_uid1054_bh793_uid1331_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1331_Out0_copy1332; -- output copy to hold a pipeline register if needed

   bh793_w80_14 <= Compressor_14_3_F200_uid1054_bh793_uid1331_Out0(0);
   bh793_w81_11 <= Compressor_14_3_F200_uid1054_bh793_uid1331_Out0(1);
   bh793_w82_11 <= Compressor_14_3_F200_uid1054_bh793_uid1331_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1333_In0 <= "" & bh793_w81_9 & bh793_w81_8 & bh793_w81_7;
   Compressor_3_2_F200_uid1040_uid1333: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1333_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1333_Out0_copy1334);
   Compressor_3_2_F200_uid1040_bh793_uid1333_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1333_Out0_copy1334; -- output copy to hold a pipeline register if needed

   bh793_w81_12 <= Compressor_3_2_F200_uid1040_bh793_uid1333_Out0(0);
   bh793_w82_12 <= Compressor_3_2_F200_uid1040_bh793_uid1333_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1335_In0 <= "" & bh793_w82_10 & bh793_w82_9 & bh793_w82_8 & bh793_w82_7;
   Compressor_14_3_F200_uid1054_bh793_uid1335_In1 <= "" & bh793_w83_9;
   Compressor_14_3_F200_uid1054_uid1335: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1335_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1335_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1335_Out0_copy1336);
   Compressor_14_3_F200_uid1054_bh793_uid1335_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1335_Out0_copy1336; -- output copy to hold a pipeline register if needed

   bh793_w82_13 <= Compressor_14_3_F200_uid1054_bh793_uid1335_Out0(0);
   bh793_w83_10 <= Compressor_14_3_F200_uid1054_bh793_uid1335_Out0(1);
   bh793_w84_9 <= Compressor_14_3_F200_uid1054_bh793_uid1335_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1337_In0 <= "" & bh793_w83_8 & bh793_w83_7 & bh793_w83_6;
   Compressor_23_3_F200_uid1032_bh793_uid1337_In1 <= "" & bh793_w84_8 & bh793_w84_7;
   Compressor_23_3_F200_uid1032_uid1337: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1337_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1337_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1337_Out0_copy1338);
   Compressor_23_3_F200_uid1032_bh793_uid1337_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1337_Out0_copy1338; -- output copy to hold a pipeline register if needed

   bh793_w83_11 <= Compressor_23_3_F200_uid1032_bh793_uid1337_Out0(0);
   bh793_w84_10 <= Compressor_23_3_F200_uid1032_bh793_uid1337_Out0(1);
   bh793_w85_10 <= Compressor_23_3_F200_uid1032_bh793_uid1337_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1339_In0 <= "" & bh793_w85_9 & bh793_w85_8 & bh793_w85_7 & bh793_w85_6;
   Compressor_14_3_F200_uid1054_bh793_uid1339_In1 <= "" & "0";
   Compressor_14_3_F200_uid1054_uid1339: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1339_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1339_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1339_Out0_copy1340);
   Compressor_14_3_F200_uid1054_bh793_uid1339_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1339_Out0_copy1340; -- output copy to hold a pipeline register if needed

   bh793_w85_11 <= Compressor_14_3_F200_uid1054_bh793_uid1339_Out0(0);
   bh793_w86_9 <= Compressor_14_3_F200_uid1054_bh793_uid1339_Out0(1);
   bh793_w87_9 <= Compressor_14_3_F200_uid1054_bh793_uid1339_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1341_In0 <= "" & bh793_w86_8 & bh793_w86_7 & bh793_w86_6;
   Compressor_3_2_F200_uid1040_uid1341: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1341_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1341_Out0_copy1342);
   Compressor_3_2_F200_uid1040_bh793_uid1341_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1341_Out0_copy1342; -- output copy to hold a pipeline register if needed

   bh793_w86_10 <= Compressor_3_2_F200_uid1040_bh793_uid1341_Out0(0);
   bh793_w87_10 <= Compressor_3_2_F200_uid1040_bh793_uid1341_Out0(1);

   Compressor_3_2_F200_uid1040_bh793_uid1343_In0 <= "" & bh793_w87_8 & bh793_w87_7 & bh793_w87_6;
   Compressor_3_2_F200_uid1040_uid1343: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1343_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1343_Out0_copy1344);
   Compressor_3_2_F200_uid1040_bh793_uid1343_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1343_Out0_copy1344; -- output copy to hold a pipeline register if needed

   bh793_w87_11 <= Compressor_3_2_F200_uid1040_bh793_uid1343_Out0(0);
   bh793_w88_10 <= Compressor_3_2_F200_uid1040_bh793_uid1343_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1345_In0 <= "" & bh793_w88_9 & bh793_w88_8 & bh793_w88_7 & bh793_w88_6;
   Compressor_14_3_F200_uid1054_bh793_uid1345_In1 <= "" & "0";
   Compressor_14_3_F200_uid1054_uid1345: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1345_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1345_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1345_Out0_copy1346);
   Compressor_14_3_F200_uid1054_bh793_uid1345_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1345_Out0_copy1346; -- output copy to hold a pipeline register if needed

   bh793_w88_11 <= Compressor_14_3_F200_uid1054_bh793_uid1345_Out0(0);
   bh793_w89_9 <= Compressor_14_3_F200_uid1054_bh793_uid1345_Out0(1);
   bh793_w90_9 <= Compressor_14_3_F200_uid1054_bh793_uid1345_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1347_In0 <= "" & bh793_w89_8 & bh793_w89_7 & bh793_w89_6;
   Compressor_3_2_F200_uid1040_uid1347: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1347_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1347_Out0_copy1348);
   Compressor_3_2_F200_uid1040_bh793_uid1347_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1347_Out0_copy1348; -- output copy to hold a pipeline register if needed

   bh793_w89_10 <= Compressor_3_2_F200_uid1040_bh793_uid1347_Out0(0);
   bh793_w90_10 <= Compressor_3_2_F200_uid1040_bh793_uid1347_Out0(1);

   Compressor_3_2_F200_uid1040_bh793_uid1349_In0 <= "" & bh793_w90_8 & bh793_w90_7 & bh793_w90_6;
   Compressor_3_2_F200_uid1040_uid1349: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1349_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1349_Out0_copy1350);
   Compressor_3_2_F200_uid1040_bh793_uid1349_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1349_Out0_copy1350; -- output copy to hold a pipeline register if needed

   bh793_w90_11 <= Compressor_3_2_F200_uid1040_bh793_uid1349_Out0(0);
   bh793_w91_10 <= Compressor_3_2_F200_uid1040_bh793_uid1349_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1351_In0 <= "" & bh793_w91_9 & bh793_w91_8 & bh793_w91_7 & bh793_w91_6;
   Compressor_14_3_F200_uid1054_bh793_uid1351_In1 <= "" & "0";
   Compressor_14_3_F200_uid1054_uid1351: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1351_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1351_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1351_Out0_copy1352);
   Compressor_14_3_F200_uid1054_bh793_uid1351_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1351_Out0_copy1352; -- output copy to hold a pipeline register if needed

   bh793_w91_11 <= Compressor_14_3_F200_uid1054_bh793_uid1351_Out0(0);
   bh793_w92_9 <= Compressor_14_3_F200_uid1054_bh793_uid1351_Out0(1);
   bh793_w93_9 <= Compressor_14_3_F200_uid1054_bh793_uid1351_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1353_In0 <= "" & bh793_w92_8 & bh793_w92_7 & bh793_w92_6;
   Compressor_3_2_F200_uid1040_uid1353: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1353_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1353_Out0_copy1354);
   Compressor_3_2_F200_uid1040_bh793_uid1353_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1353_Out0_copy1354; -- output copy to hold a pipeline register if needed

   bh793_w92_10 <= Compressor_3_2_F200_uid1040_bh793_uid1353_Out0(0);
   bh793_w93_10 <= Compressor_3_2_F200_uid1040_bh793_uid1353_Out0(1);

   Compressor_3_2_F200_uid1040_bh793_uid1355_In0 <= "" & bh793_w93_8 & bh793_w93_7 & bh793_w93_6;
   Compressor_3_2_F200_uid1040_uid1355: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1355_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1355_Out0_copy1356);
   Compressor_3_2_F200_uid1040_bh793_uid1355_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1355_Out0_copy1356; -- output copy to hold a pipeline register if needed

   bh793_w93_11 <= Compressor_3_2_F200_uid1040_bh793_uid1355_Out0(0);
   bh793_w94_10 <= Compressor_3_2_F200_uid1040_bh793_uid1355_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1357_In0 <= "" & bh793_w94_9 & bh793_w94_8 & bh793_w94_7 & bh793_w94_6;
   Compressor_14_3_F200_uid1054_bh793_uid1357_In1 <= "" & "0";
   Compressor_14_3_F200_uid1054_uid1357: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1357_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1357_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1357_Out0_copy1358);
   Compressor_14_3_F200_uid1054_bh793_uid1357_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1357_Out0_copy1358; -- output copy to hold a pipeline register if needed

   bh793_w94_11 <= Compressor_14_3_F200_uid1054_bh793_uid1357_Out0(0);
   bh793_w95_9 <= Compressor_14_3_F200_uid1054_bh793_uid1357_Out0(1);
   bh793_w96_9 <= Compressor_14_3_F200_uid1054_bh793_uid1357_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1359_In0 <= "" & bh793_w95_8 & bh793_w95_7 & bh793_w95_6;
   Compressor_3_2_F200_uid1040_uid1359: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1359_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1359_Out0_copy1360);
   Compressor_3_2_F200_uid1040_bh793_uid1359_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1359_Out0_copy1360; -- output copy to hold a pipeline register if needed

   bh793_w95_10 <= Compressor_3_2_F200_uid1040_bh793_uid1359_Out0(0);
   bh793_w96_10 <= Compressor_3_2_F200_uid1040_bh793_uid1359_Out0(1);

   Compressor_3_2_F200_uid1040_bh793_uid1361_In0 <= "" & bh793_w96_8 & bh793_w96_7 & bh793_w96_6;
   Compressor_3_2_F200_uid1040_uid1361: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1361_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1361_Out0_copy1362);
   Compressor_3_2_F200_uid1040_bh793_uid1361_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1361_Out0_copy1362; -- output copy to hold a pipeline register if needed

   bh793_w96_11 <= Compressor_3_2_F200_uid1040_bh793_uid1361_Out0(0);
   bh793_w97_10 <= Compressor_3_2_F200_uid1040_bh793_uid1361_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1363_In0 <= "" & bh793_w97_9 & bh793_w97_8 & bh793_w97_7 & bh793_w97_6;
   Compressor_14_3_F200_uid1054_bh793_uid1363_In1 <= "" & "0";
   Compressor_14_3_F200_uid1054_uid1363: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1363_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1363_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1363_Out0_copy1364);
   Compressor_14_3_F200_uid1054_bh793_uid1363_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1363_Out0_copy1364; -- output copy to hold a pipeline register if needed

   bh793_w97_11 <= Compressor_14_3_F200_uid1054_bh793_uid1363_Out0(0);
   bh793_w98_9 <= Compressor_14_3_F200_uid1054_bh793_uid1363_Out0(1);
   bh793_w99_9 <= Compressor_14_3_F200_uid1054_bh793_uid1363_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1365_In0 <= "" & bh793_w98_8 & bh793_w98_7 & bh793_w98_6;
   Compressor_3_2_F200_uid1040_uid1365: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1365_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1365_Out0_copy1366);
   Compressor_3_2_F200_uid1040_bh793_uid1365_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1365_Out0_copy1366; -- output copy to hold a pipeline register if needed

   bh793_w98_10 <= Compressor_3_2_F200_uid1040_bh793_uid1365_Out0(0);
   bh793_w99_10 <= Compressor_3_2_F200_uid1040_bh793_uid1365_Out0(1);

   Compressor_23_3_F200_uid1032_bh793_uid1367_In0 <= "" & bh793_w99_8 & bh793_w99_7 & bh793_w99_6;
   Compressor_23_3_F200_uid1032_bh793_uid1367_In1 <= "" & bh793_w100_8 & bh793_w100_7;
   Compressor_23_3_F200_uid1032_uid1367: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1367_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1367_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1367_Out0_copy1368);
   Compressor_23_3_F200_uid1032_bh793_uid1367_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1367_Out0_copy1368; -- output copy to hold a pipeline register if needed

   bh793_w99_11 <= Compressor_23_3_F200_uid1032_bh793_uid1367_Out0(0);
   bh793_w100_9 <= Compressor_23_3_F200_uid1032_bh793_uid1367_Out0(1);
   bh793_w101_6 <= Compressor_23_3_F200_uid1032_bh793_uid1367_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1369_In0 <= "" & bh793_w101_5 & bh793_w101_4 & bh793_w101_3;
   Compressor_23_3_F200_uid1032_bh793_uid1369_In1 <= "" & bh793_w102_6 & bh793_w102_5;
   Compressor_23_3_F200_uid1032_uid1369: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1369_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1369_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1369_Out0_copy1370);
   Compressor_23_3_F200_uid1032_bh793_uid1369_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1369_Out0_copy1370; -- output copy to hold a pipeline register if needed

   bh793_w101_7 <= Compressor_23_3_F200_uid1032_bh793_uid1369_Out0(0);
   bh793_w102_7 <= Compressor_23_3_F200_uid1032_bh793_uid1369_Out0(1);
   bh793_w103_3 <= Compressor_23_3_F200_uid1032_bh793_uid1369_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1371_In0 <= "" & bh793_w103_2 & bh793_w103_1 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1371_In1 <= "" & bh793_w104_1 & bh793_w104_0;
   Compressor_23_3_F200_uid1032_uid1371: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1371_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1371_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1371_Out0_copy1372);
   Compressor_23_3_F200_uid1032_bh793_uid1371_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1371_Out0_copy1372; -- output copy to hold a pipeline register if needed

   bh793_w103_4 <= Compressor_23_3_F200_uid1032_bh793_uid1371_Out0(0);
   bh793_w104_2 <= Compressor_23_3_F200_uid1032_bh793_uid1371_Out0(1);
   bh793_w105_1 <= Compressor_23_3_F200_uid1032_bh793_uid1371_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1373_In0 <= "" & bh793_w21_5 & bh793_w21_4 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1373_In1 <= "" & bh793_w22_3;
   Compressor_14_3_F200_uid1054_uid1373: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1373_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1373_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1373_Out0_copy1374);
   Compressor_14_3_F200_uid1054_bh793_uid1373_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1373_Out0_copy1374; -- output copy to hold a pipeline register if needed

   bh793_w21_6 <= Compressor_14_3_F200_uid1054_bh793_uid1373_Out0(0);
   bh793_w22_4 <= Compressor_14_3_F200_uid1054_bh793_uid1373_Out0(1);
   bh793_w23_6 <= Compressor_14_3_F200_uid1054_bh793_uid1373_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1375_In0 <= "" & bh793_w23_5 & bh793_w23_4 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1375_In1 <= "" & bh793_w24_5;
   Compressor_14_3_F200_uid1054_uid1375: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1375_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1375_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1375_Out0_copy1376);
   Compressor_14_3_F200_uid1054_bh793_uid1375_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1375_Out0_copy1376; -- output copy to hold a pipeline register if needed

   bh793_w23_7 <= Compressor_14_3_F200_uid1054_bh793_uid1375_Out0(0);
   bh793_w24_6 <= Compressor_14_3_F200_uid1054_bh793_uid1375_Out0(1);
   bh793_w25_6 <= Compressor_14_3_F200_uid1054_bh793_uid1375_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1377_In0 <= "" & bh793_w25_5 & bh793_w25_4 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1377_In1 <= "" & bh793_w26_5;
   Compressor_14_3_F200_uid1054_uid1377: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1377_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1377_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1377_Out0_copy1378);
   Compressor_14_3_F200_uid1054_bh793_uid1377_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1377_Out0_copy1378; -- output copy to hold a pipeline register if needed

   bh793_w25_7 <= Compressor_14_3_F200_uid1054_bh793_uid1377_Out0(0);
   bh793_w26_6 <= Compressor_14_3_F200_uid1054_bh793_uid1377_Out0(1);
   bh793_w27_6 <= Compressor_14_3_F200_uid1054_bh793_uid1377_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1379_In0 <= "" & bh793_w27_5 & bh793_w27_4 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1379_In1 <= "" & bh793_w28_5;
   Compressor_14_3_F200_uid1054_uid1379: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1379_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1379_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1379_Out0_copy1380);
   Compressor_14_3_F200_uid1054_bh793_uid1379_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1379_Out0_copy1380; -- output copy to hold a pipeline register if needed

   bh793_w27_7 <= Compressor_14_3_F200_uid1054_bh793_uid1379_Out0(0);
   bh793_w28_6 <= Compressor_14_3_F200_uid1054_bh793_uid1379_Out0(1);
   bh793_w29_6 <= Compressor_14_3_F200_uid1054_bh793_uid1379_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1381_In0 <= "" & bh793_w29_5 & bh793_w29_4 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1381_In1 <= "" & bh793_w30_5;
   Compressor_14_3_F200_uid1054_uid1381: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1381_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1381_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1381_Out0_copy1382);
   Compressor_14_3_F200_uid1054_bh793_uid1381_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1381_Out0_copy1382; -- output copy to hold a pipeline register if needed

   bh793_w29_7 <= Compressor_14_3_F200_uid1054_bh793_uid1381_Out0(0);
   bh793_w30_6 <= Compressor_14_3_F200_uid1054_bh793_uid1381_Out0(1);
   bh793_w31_6 <= Compressor_14_3_F200_uid1054_bh793_uid1381_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1383_In0 <= "" & bh793_w31_5 & bh793_w31_4 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1383_In1 <= "" & bh793_w32_5;
   Compressor_14_3_F200_uid1054_uid1383: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1383_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1383_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1383_Out0_copy1384);
   Compressor_14_3_F200_uid1054_bh793_uid1383_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1383_Out0_copy1384; -- output copy to hold a pipeline register if needed

   bh793_w31_7 <= Compressor_14_3_F200_uid1054_bh793_uid1383_Out0(0);
   bh793_w32_6 <= Compressor_14_3_F200_uid1054_bh793_uid1383_Out0(1);
   bh793_w33_6 <= Compressor_14_3_F200_uid1054_bh793_uid1383_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1385_In0 <= "" & bh793_w33_5 & bh793_w33_4 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1385_In1 <= "" & bh793_w34_6;
   Compressor_14_3_F200_uid1054_uid1385: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1385_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1385_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1385_Out0_copy1386);
   Compressor_14_3_F200_uid1054_bh793_uid1385_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1385_Out0_copy1386; -- output copy to hold a pipeline register if needed

   bh793_w33_7 <= Compressor_14_3_F200_uid1054_bh793_uid1385_Out0(0);
   bh793_w34_7 <= Compressor_14_3_F200_uid1054_bh793_uid1385_Out0(1);
   bh793_w35_8 <= Compressor_14_3_F200_uid1054_bh793_uid1385_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1387_In0 <= "" & bh793_w35_7 & bh793_w35_6 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1387_In1 <= "" & bh793_w36_8 & bh793_w36_7;
   Compressor_23_3_F200_uid1032_uid1387: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1387_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1387_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1387_Out0_copy1388);
   Compressor_23_3_F200_uid1032_bh793_uid1387_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1387_Out0_copy1388; -- output copy to hold a pipeline register if needed

   bh793_w35_9 <= Compressor_23_3_F200_uid1032_bh793_uid1387_Out0(0);
   bh793_w36_9 <= Compressor_23_3_F200_uid1032_bh793_uid1387_Out0(1);
   bh793_w37_7 <= Compressor_23_3_F200_uid1032_bh793_uid1387_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1389_In0 <= "" & bh793_w38_8 & bh793_w38_7 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1389_In1 <= "" & bh793_w39_6;
   Compressor_14_3_F200_uid1054_uid1389: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1389_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1389_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1389_Out0_copy1390);
   Compressor_14_3_F200_uid1054_bh793_uid1389_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1389_Out0_copy1390; -- output copy to hold a pipeline register if needed

   bh793_w38_9 <= Compressor_14_3_F200_uid1054_bh793_uid1389_Out0(0);
   bh793_w39_7 <= Compressor_14_3_F200_uid1054_bh793_uid1389_Out0(1);
   bh793_w40_9 <= Compressor_14_3_F200_uid1054_bh793_uid1389_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1391_In0 <= "" & bh793_w40_8 & bh793_w40_7 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1391_In1 <= "" & bh793_w41_6;
   Compressor_14_3_F200_uid1054_uid1391: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1391_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1391_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1391_Out0_copy1392);
   Compressor_14_3_F200_uid1054_bh793_uid1391_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1391_Out0_copy1392; -- output copy to hold a pipeline register if needed

   bh793_w40_10 <= Compressor_14_3_F200_uid1054_bh793_uid1391_Out0(0);
   bh793_w41_7 <= Compressor_14_3_F200_uid1054_bh793_uid1391_Out0(1);
   bh793_w42_9 <= Compressor_14_3_F200_uid1054_bh793_uid1391_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1393_In0 <= "" & bh793_w42_8 & bh793_w42_7 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1393_In1 <= "" & bh793_w43_6;
   Compressor_14_3_F200_uid1054_uid1393: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1393_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1393_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1393_Out0_copy1394);
   Compressor_14_3_F200_uid1054_bh793_uid1393_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1393_Out0_copy1394; -- output copy to hold a pipeline register if needed

   bh793_w42_10 <= Compressor_14_3_F200_uid1054_bh793_uid1393_Out0(0);
   bh793_w43_7 <= Compressor_14_3_F200_uid1054_bh793_uid1393_Out0(1);
   bh793_w44_9 <= Compressor_14_3_F200_uid1054_bh793_uid1393_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1395_In0 <= "" & bh793_w44_8 & bh793_w44_7 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1395_In1 <= "" & bh793_w45_6;
   Compressor_14_3_F200_uid1054_uid1395: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1395_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1395_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1395_Out0_copy1396);
   Compressor_14_3_F200_uid1054_bh793_uid1395_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1395_Out0_copy1396; -- output copy to hold a pipeline register if needed

   bh793_w44_10 <= Compressor_14_3_F200_uid1054_bh793_uid1395_Out0(0);
   bh793_w45_7 <= Compressor_14_3_F200_uid1054_bh793_uid1395_Out0(1);
   bh793_w46_9 <= Compressor_14_3_F200_uid1054_bh793_uid1395_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1397_In0 <= "" & bh793_w46_8 & bh793_w46_7 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1397_In1 <= "" & bh793_w47_6;
   Compressor_14_3_F200_uid1054_uid1397: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1397_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1397_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1397_Out0_copy1398);
   Compressor_14_3_F200_uid1054_bh793_uid1397_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1397_Out0_copy1398; -- output copy to hold a pipeline register if needed

   bh793_w46_10 <= Compressor_14_3_F200_uid1054_bh793_uid1397_Out0(0);
   bh793_w47_7 <= Compressor_14_3_F200_uid1054_bh793_uid1397_Out0(1);
   bh793_w48_10 <= Compressor_14_3_F200_uid1054_bh793_uid1397_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1399_In0 <= "" & bh793_w48_9 & bh793_w48_8 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1399_In1 <= "" & bh793_w49_7 & bh793_w49_8;
   Compressor_23_3_F200_uid1032_uid1399: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1399_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1399_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1399_Out0_copy1400);
   Compressor_23_3_F200_uid1032_bh793_uid1399_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1399_Out0_copy1400; -- output copy to hold a pipeline register if needed

   bh793_w48_11 <= Compressor_23_3_F200_uid1032_bh793_uid1399_Out0(0);
   bh793_w49_9 <= Compressor_23_3_F200_uid1032_bh793_uid1399_Out0(1);
   bh793_w50_12 <= Compressor_23_3_F200_uid1032_bh793_uid1399_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1401_In0 <= "" & bh793_w50_9 & bh793_w50_11 & bh793_w50_10;
   Compressor_23_3_F200_uid1032_bh793_uid1401_In1 <= "" & bh793_w51_11 & bh793_w51_8;
   Compressor_23_3_F200_uid1032_uid1401: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1401_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1401_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1401_Out0_copy1402);
   Compressor_23_3_F200_uid1032_bh793_uid1401_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1401_Out0_copy1402; -- output copy to hold a pipeline register if needed

   bh793_w50_13 <= Compressor_23_3_F200_uid1032_bh793_uid1401_Out0(0);
   bh793_w51_12 <= Compressor_23_3_F200_uid1032_bh793_uid1401_Out0(1);
   bh793_w52_16 <= Compressor_23_3_F200_uid1032_bh793_uid1401_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1403_In0 <= "" & bh793_w52_15 & bh793_w52_14 & bh793_w52_9;
   Compressor_23_3_F200_uid1032_bh793_uid1403_In1 <= "" & bh793_w53_14 & bh793_w53_13;
   Compressor_23_3_F200_uid1032_uid1403: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1403_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1403_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1403_Out0_copy1404);
   Compressor_23_3_F200_uid1032_bh793_uid1403_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1403_Out0_copy1404; -- output copy to hold a pipeline register if needed

   bh793_w52_17 <= Compressor_23_3_F200_uid1032_bh793_uid1403_Out0(0);
   bh793_w53_15 <= Compressor_23_3_F200_uid1032_bh793_uid1403_Out0(1);
   bh793_w54_18 <= Compressor_23_3_F200_uid1032_bh793_uid1403_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1405_In0 <= "" & bh793_w54_16 & bh793_w54_17 & bh793_w54_15;
   Compressor_3_2_F200_uid1040_uid1405: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1405_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1405_Out0_copy1406);
   Compressor_3_2_F200_uid1040_bh793_uid1405_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1405_Out0_copy1406; -- output copy to hold a pipeline register if needed

   bh793_w54_19 <= Compressor_3_2_F200_uid1040_bh793_uid1405_Out0(0);
   bh793_w55_17 <= Compressor_3_2_F200_uid1040_bh793_uid1405_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1407_In0 <= "" & bh793_w55_14 & bh793_w55_15 & bh793_w55_16 & bh793_w55_9;
   Compressor_14_3_F200_uid1054_bh793_uid1407_In1 <= "" & "0";
   Compressor_14_3_F200_uid1054_uid1407: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1407_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1407_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1407_Out0_copy1408);
   Compressor_14_3_F200_uid1054_bh793_uid1407_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1407_Out0_copy1408; -- output copy to hold a pipeline register if needed

   bh793_w55_18 <= Compressor_14_3_F200_uid1054_bh793_uid1407_Out0(0);
   bh793_w56_18 <= Compressor_14_3_F200_uid1054_bh793_uid1407_Out0(1);
   bh793_w57_17 <= Compressor_14_3_F200_uid1054_bh793_uid1407_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1409_In0 <= "" & bh793_w56_15 & bh793_w56_17 & bh793_w56_16;
   Compressor_3_2_F200_uid1040_uid1409: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1409_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1409_Out0_copy1410);
   Compressor_3_2_F200_uid1040_bh793_uid1409_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1409_Out0_copy1410; -- output copy to hold a pipeline register if needed

   bh793_w56_19 <= Compressor_3_2_F200_uid1040_bh793_uid1409_Out0(0);
   bh793_w57_18 <= Compressor_3_2_F200_uid1040_bh793_uid1409_Out0(1);

   Compressor_3_2_F200_uid1040_bh793_uid1411_In0 <= "" & bh793_w57_15 & bh793_w57_16 & bh793_w57_10;
   Compressor_3_2_F200_uid1040_uid1411: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1411_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1411_Out0_copy1412);
   Compressor_3_2_F200_uid1040_bh793_uid1411_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1411_Out0_copy1412; -- output copy to hold a pipeline register if needed

   bh793_w57_19 <= Compressor_3_2_F200_uid1040_bh793_uid1411_Out0(0);
   bh793_w58_17 <= Compressor_3_2_F200_uid1040_bh793_uid1411_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1413_In0 <= "" & bh793_w58_14 & bh793_w58_15 & bh793_w58_16 & bh793_w58_9;
   Compressor_14_3_F200_uid1054_bh793_uid1413_In1 <= "" & "0";
   Compressor_14_3_F200_uid1054_uid1413: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1413_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1413_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1413_Out0_copy1414);
   Compressor_14_3_F200_uid1054_bh793_uid1413_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1413_Out0_copy1414; -- output copy to hold a pipeline register if needed

   bh793_w58_18 <= Compressor_14_3_F200_uid1054_bh793_uid1413_Out0(0);
   bh793_w59_18 <= Compressor_14_3_F200_uid1054_bh793_uid1413_Out0(1);
   bh793_w60_17 <= Compressor_14_3_F200_uid1054_bh793_uid1413_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1415_In0 <= "" & bh793_w59_15 & bh793_w59_17 & bh793_w59_16;
   Compressor_3_2_F200_uid1040_uid1415: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1415_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1415_Out0_copy1416);
   Compressor_3_2_F200_uid1040_bh793_uid1415_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1415_Out0_copy1416; -- output copy to hold a pipeline register if needed

   bh793_w59_19 <= Compressor_3_2_F200_uid1040_bh793_uid1415_Out0(0);
   bh793_w60_18 <= Compressor_3_2_F200_uid1040_bh793_uid1415_Out0(1);

   Compressor_3_2_F200_uid1040_bh793_uid1417_In0 <= "" & bh793_w60_15 & bh793_w60_16 & bh793_w60_10;
   Compressor_3_2_F200_uid1040_uid1417: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1417_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1417_Out0_copy1418);
   Compressor_3_2_F200_uid1040_bh793_uid1417_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1417_Out0_copy1418; -- output copy to hold a pipeline register if needed

   bh793_w60_19 <= Compressor_3_2_F200_uid1040_bh793_uid1417_Out0(0);
   bh793_w61_17 <= Compressor_3_2_F200_uid1040_bh793_uid1417_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1419_In0 <= "" & bh793_w61_14 & bh793_w61_15 & bh793_w61_16 & bh793_w61_9;
   Compressor_14_3_F200_uid1054_bh793_uid1419_In1 <= "" & "0";
   Compressor_14_3_F200_uid1054_uid1419: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1419_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1419_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1419_Out0_copy1420);
   Compressor_14_3_F200_uid1054_bh793_uid1419_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1419_Out0_copy1420; -- output copy to hold a pipeline register if needed

   bh793_w61_18 <= Compressor_14_3_F200_uid1054_bh793_uid1419_Out0(0);
   bh793_w62_18 <= Compressor_14_3_F200_uid1054_bh793_uid1419_Out0(1);
   bh793_w63_17 <= Compressor_14_3_F200_uid1054_bh793_uid1419_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1421_In0 <= "" & bh793_w62_15 & bh793_w62_17 & bh793_w62_16;
   Compressor_3_2_F200_uid1040_uid1421: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1421_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1421_Out0_copy1422);
   Compressor_3_2_F200_uid1040_bh793_uid1421_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1421_Out0_copy1422; -- output copy to hold a pipeline register if needed

   bh793_w62_19 <= Compressor_3_2_F200_uid1040_bh793_uid1421_Out0(0);
   bh793_w63_18 <= Compressor_3_2_F200_uid1040_bh793_uid1421_Out0(1);

   Compressor_3_2_F200_uid1040_bh793_uid1423_In0 <= "" & bh793_w63_15 & bh793_w63_16 & bh793_w63_10;
   Compressor_3_2_F200_uid1040_uid1423: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1423_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1423_Out0_copy1424);
   Compressor_3_2_F200_uid1040_bh793_uid1423_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1423_Out0_copy1424; -- output copy to hold a pipeline register if needed

   bh793_w63_19 <= Compressor_3_2_F200_uid1040_bh793_uid1423_Out0(0);
   bh793_w64_17 <= Compressor_3_2_F200_uid1040_bh793_uid1423_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1425_In0 <= "" & bh793_w64_14 & bh793_w64_15 & bh793_w64_16 & bh793_w64_9;
   Compressor_14_3_F200_uid1054_bh793_uid1425_In1 <= "" & "0";
   Compressor_14_3_F200_uid1054_uid1425: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1425_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1425_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1425_Out0_copy1426);
   Compressor_14_3_F200_uid1054_bh793_uid1425_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1425_Out0_copy1426; -- output copy to hold a pipeline register if needed

   bh793_w64_18 <= Compressor_14_3_F200_uid1054_bh793_uid1425_Out0(0);
   bh793_w65_18 <= Compressor_14_3_F200_uid1054_bh793_uid1425_Out0(1);
   bh793_w66_16 <= Compressor_14_3_F200_uid1054_bh793_uid1425_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1427_In0 <= "" & bh793_w65_15 & bh793_w65_17 & bh793_w65_16;
   Compressor_3_2_F200_uid1040_uid1427: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1427_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1427_Out0_copy1428);
   Compressor_3_2_F200_uid1040_bh793_uid1427_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1427_Out0_copy1428; -- output copy to hold a pipeline register if needed

   bh793_w65_19 <= Compressor_3_2_F200_uid1040_bh793_uid1427_Out0(0);
   bh793_w66_17 <= Compressor_3_2_F200_uid1040_bh793_uid1427_Out0(1);

   Compressor_23_3_F200_uid1032_bh793_uid1429_In0 <= "" & bh793_w66_14 & bh793_w66_15 & bh793_w66_9;
   Compressor_23_3_F200_uid1032_bh793_uid1429_In1 <= "" & bh793_w67_13 & bh793_w67_14;
   Compressor_23_3_F200_uid1032_uid1429: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1429_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1429_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1429_Out0_copy1430);
   Compressor_23_3_F200_uid1032_bh793_uid1429_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1429_Out0_copy1430; -- output copy to hold a pipeline register if needed

   bh793_w66_18 <= Compressor_23_3_F200_uid1032_bh793_uid1429_Out0(0);
   bh793_w67_16 <= Compressor_23_3_F200_uid1032_bh793_uid1429_Out0(1);
   bh793_w68_17 <= Compressor_23_3_F200_uid1032_bh793_uid1429_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1431_In0 <= "" & bh793_w68_14 & bh793_w68_16 & bh793_w68_15;
   Compressor_23_3_F200_uid1032_bh793_uid1431_In1 <= "" & bh793_w69_14 & bh793_w69_13;
   Compressor_23_3_F200_uid1032_uid1431: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1431_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1431_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1431_Out0_copy1432);
   Compressor_23_3_F200_uid1032_bh793_uid1431_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1431_Out0_copy1432; -- output copy to hold a pipeline register if needed

   bh793_w68_18 <= Compressor_23_3_F200_uid1032_bh793_uid1431_Out0(0);
   bh793_w69_15 <= Compressor_23_3_F200_uid1032_bh793_uid1431_Out0(1);
   bh793_w70_16 <= Compressor_23_3_F200_uid1032_bh793_uid1431_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1433_In0 <= "" & bh793_w70_15 & bh793_w70_14 & bh793_w70_13 & bh793_w70_8;
   Compressor_14_3_F200_uid1054_bh793_uid1433_In1 <= "" & bh793_w71_15;
   Compressor_14_3_F200_uid1054_uid1433: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1433_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1433_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1433_Out0_copy1434);
   Compressor_14_3_F200_uid1054_bh793_uid1433_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1433_Out0_copy1434; -- output copy to hold a pipeline register if needed

   bh793_w70_17 <= Compressor_14_3_F200_uid1054_bh793_uid1433_Out0(0);
   bh793_w71_16 <= Compressor_14_3_F200_uid1054_bh793_uid1433_Out0(1);
   bh793_w72_15 <= Compressor_14_3_F200_uid1054_bh793_uid1433_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1435_In0 <= "" & bh793_w72_14 & bh793_w72_13 & bh793_w72_12;
   Compressor_3_2_F200_uid1040_uid1435: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1435_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1435_Out0_copy1436);
   Compressor_3_2_F200_uid1040_bh793_uid1435_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1435_Out0_copy1436; -- output copy to hold a pipeline register if needed

   bh793_w72_16 <= Compressor_3_2_F200_uid1040_bh793_uid1435_Out0(0);
   bh793_w73_16 <= Compressor_3_2_F200_uid1040_bh793_uid1435_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1437_In0 <= "" & bh793_w73_15 & bh793_w73_14 & bh793_w73_13 & bh793_w73_8;
   Compressor_14_3_F200_uid1054_bh793_uid1437_In1 <= "" & bh793_w74_15;
   Compressor_14_3_F200_uid1054_uid1437: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1437_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1437_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1437_Out0_copy1438);
   Compressor_14_3_F200_uid1054_bh793_uid1437_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1437_Out0_copy1438; -- output copy to hold a pipeline register if needed

   bh793_w73_17 <= Compressor_14_3_F200_uid1054_bh793_uid1437_Out0(0);
   bh793_w74_16 <= Compressor_14_3_F200_uid1054_bh793_uid1437_Out0(1);
   bh793_w75_15 <= Compressor_14_3_F200_uid1054_bh793_uid1437_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1439_In0 <= "" & bh793_w75_14 & bh793_w75_13 & bh793_w75_12;
   Compressor_3_2_F200_uid1040_uid1439: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1439_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1439_Out0_copy1440);
   Compressor_3_2_F200_uid1040_bh793_uid1439_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1439_Out0_copy1440; -- output copy to hold a pipeline register if needed

   bh793_w75_16 <= Compressor_3_2_F200_uid1040_bh793_uid1439_Out0(0);
   bh793_w76_16 <= Compressor_3_2_F200_uid1040_bh793_uid1439_Out0(1);

   Compressor_14_3_F200_uid1054_bh793_uid1441_In0 <= "" & bh793_w76_15 & bh793_w76_14 & bh793_w76_13 & bh793_w76_8;
   Compressor_14_3_F200_uid1054_bh793_uid1441_In1 <= "" & bh793_w77_13;
   Compressor_14_3_F200_uid1054_uid1441: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1441_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1441_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1441_Out0_copy1442);
   Compressor_14_3_F200_uid1054_bh793_uid1441_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1441_Out0_copy1442; -- output copy to hold a pipeline register if needed

   bh793_w76_17 <= Compressor_14_3_F200_uid1054_bh793_uid1441_Out0(0);
   bh793_w77_14 <= Compressor_14_3_F200_uid1054_bh793_uid1441_Out0(1);
   bh793_w78_14 <= Compressor_14_3_F200_uid1054_bh793_uid1441_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1443_In0 <= "" & bh793_w78_13 & bh793_w78_12 & bh793_w78_11 & bh793_w78_6;
   Compressor_14_3_F200_uid1054_bh793_uid1443_In1 <= "" & bh793_w79_11;
   Compressor_14_3_F200_uid1054_uid1443: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1443_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1443_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1443_Out0_copy1444);
   Compressor_14_3_F200_uid1054_bh793_uid1443_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1443_Out0_copy1444; -- output copy to hold a pipeline register if needed

   bh793_w78_15 <= Compressor_14_3_F200_uid1054_bh793_uid1443_Out0(0);
   bh793_w79_12 <= Compressor_14_3_F200_uid1054_bh793_uid1443_Out0(1);
   bh793_w80_15 <= Compressor_14_3_F200_uid1054_bh793_uid1443_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1445_In0 <= "" & bh793_w80_14 & bh793_w80_13 & bh793_w80_12;
   Compressor_23_3_F200_uid1032_bh793_uid1445_In1 <= "" & bh793_w81_12 & bh793_w81_11;
   Compressor_23_3_F200_uid1032_uid1445: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1445_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1445_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1445_Out0_copy1446);
   Compressor_23_3_F200_uid1032_bh793_uid1445_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1445_Out0_copy1446; -- output copy to hold a pipeline register if needed

   bh793_w80_16 <= Compressor_23_3_F200_uid1032_bh793_uid1445_Out0(0);
   bh793_w81_13 <= Compressor_23_3_F200_uid1032_bh793_uid1445_Out0(1);
   bh793_w82_14 <= Compressor_23_3_F200_uid1032_bh793_uid1445_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1447_In0 <= "" & bh793_w82_13 & bh793_w82_12 & bh793_w82_11 & bh793_w82_6;
   Compressor_14_3_F200_uid1054_bh793_uid1447_In1 <= "" & bh793_w83_11;
   Compressor_14_3_F200_uid1054_uid1447: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1447_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1447_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1447_Out0_copy1448);
   Compressor_14_3_F200_uid1054_bh793_uid1447_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1447_Out0_copy1448; -- output copy to hold a pipeline register if needed

   bh793_w82_15 <= Compressor_14_3_F200_uid1054_bh793_uid1447_Out0(0);
   bh793_w83_12 <= Compressor_14_3_F200_uid1054_bh793_uid1447_Out0(1);
   bh793_w84_11 <= Compressor_14_3_F200_uid1054_bh793_uid1447_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1449_In0 <= "" & bh793_w84_10 & bh793_w84_9 & bh793_w84_6;
   Compressor_23_3_F200_uid1032_bh793_uid1449_In1 <= "" & bh793_w85_11 & bh793_w85_10;
   Compressor_23_3_F200_uid1032_uid1449: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1449_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1449_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1449_Out0_copy1450);
   Compressor_23_3_F200_uid1032_bh793_uid1449_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1449_Out0_copy1450; -- output copy to hold a pipeline register if needed

   bh793_w84_12 <= Compressor_23_3_F200_uid1032_bh793_uid1449_Out0(0);
   bh793_w85_12 <= Compressor_23_3_F200_uid1032_bh793_uid1449_Out0(1);
   bh793_w86_11 <= Compressor_23_3_F200_uid1032_bh793_uid1449_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1451_In0 <= "" & bh793_w86_9 & bh793_w86_10 & "0";
   Compressor_3_2_F200_uid1040_uid1451: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1451_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1451_Out0_copy1452);
   Compressor_3_2_F200_uid1040_bh793_uid1451_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1451_Out0_copy1452; -- output copy to hold a pipeline register if needed

   bh793_w86_12 <= Compressor_3_2_F200_uid1040_bh793_uid1451_Out0(0);
   bh793_w87_12 <= Compressor_3_2_F200_uid1040_bh793_uid1451_Out0(1);

   Compressor_23_3_F200_uid1032_bh793_uid1453_In0 <= "" & bh793_w87_9 & bh793_w87_11 & bh793_w87_10;
   Compressor_23_3_F200_uid1032_bh793_uid1453_In1 <= "" & bh793_w88_11 & bh793_w88_10;
   Compressor_23_3_F200_uid1032_uid1453: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1453_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1453_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1453_Out0_copy1454);
   Compressor_23_3_F200_uid1032_bh793_uid1453_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1453_Out0_copy1454; -- output copy to hold a pipeline register if needed

   bh793_w87_13 <= Compressor_23_3_F200_uid1032_bh793_uid1453_Out0(0);
   bh793_w88_12 <= Compressor_23_3_F200_uid1032_bh793_uid1453_Out0(1);
   bh793_w89_11 <= Compressor_23_3_F200_uid1032_bh793_uid1453_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1455_In0 <= "" & bh793_w89_9 & bh793_w89_10 & "0";
   Compressor_3_2_F200_uid1040_uid1455: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1455_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1455_Out0_copy1456);
   Compressor_3_2_F200_uid1040_bh793_uid1455_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1455_Out0_copy1456; -- output copy to hold a pipeline register if needed

   bh793_w89_12 <= Compressor_3_2_F200_uid1040_bh793_uid1455_Out0(0);
   bh793_w90_12 <= Compressor_3_2_F200_uid1040_bh793_uid1455_Out0(1);

   Compressor_23_3_F200_uid1032_bh793_uid1457_In0 <= "" & bh793_w90_9 & bh793_w90_11 & bh793_w90_10;
   Compressor_23_3_F200_uid1032_bh793_uid1457_In1 <= "" & bh793_w91_11 & bh793_w91_10;
   Compressor_23_3_F200_uid1032_uid1457: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1457_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1457_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1457_Out0_copy1458);
   Compressor_23_3_F200_uid1032_bh793_uid1457_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1457_Out0_copy1458; -- output copy to hold a pipeline register if needed

   bh793_w90_13 <= Compressor_23_3_F200_uid1032_bh793_uid1457_Out0(0);
   bh793_w91_12 <= Compressor_23_3_F200_uid1032_bh793_uid1457_Out0(1);
   bh793_w92_11 <= Compressor_23_3_F200_uid1032_bh793_uid1457_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1459_In0 <= "" & bh793_w92_9 & bh793_w92_10 & "0";
   Compressor_3_2_F200_uid1040_uid1459: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1459_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1459_Out0_copy1460);
   Compressor_3_2_F200_uid1040_bh793_uid1459_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1459_Out0_copy1460; -- output copy to hold a pipeline register if needed

   bh793_w92_12 <= Compressor_3_2_F200_uid1040_bh793_uid1459_Out0(0);
   bh793_w93_12 <= Compressor_3_2_F200_uid1040_bh793_uid1459_Out0(1);

   Compressor_23_3_F200_uid1032_bh793_uid1461_In0 <= "" & bh793_w93_9 & bh793_w93_11 & bh793_w93_10;
   Compressor_23_3_F200_uid1032_bh793_uid1461_In1 <= "" & bh793_w94_11 & bh793_w94_10;
   Compressor_23_3_F200_uid1032_uid1461: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1461_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1461_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1461_Out0_copy1462);
   Compressor_23_3_F200_uid1032_bh793_uid1461_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1461_Out0_copy1462; -- output copy to hold a pipeline register if needed

   bh793_w93_13 <= Compressor_23_3_F200_uid1032_bh793_uid1461_Out0(0);
   bh793_w94_12 <= Compressor_23_3_F200_uid1032_bh793_uid1461_Out0(1);
   bh793_w95_11 <= Compressor_23_3_F200_uid1032_bh793_uid1461_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1463_In0 <= "" & bh793_w95_9 & bh793_w95_10 & "0";
   Compressor_3_2_F200_uid1040_uid1463: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1463_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1463_Out0_copy1464);
   Compressor_3_2_F200_uid1040_bh793_uid1463_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1463_Out0_copy1464; -- output copy to hold a pipeline register if needed

   bh793_w95_12 <= Compressor_3_2_F200_uid1040_bh793_uid1463_Out0(0);
   bh793_w96_12 <= Compressor_3_2_F200_uid1040_bh793_uid1463_Out0(1);

   Compressor_23_3_F200_uid1032_bh793_uid1465_In0 <= "" & bh793_w96_9 & bh793_w96_11 & bh793_w96_10;
   Compressor_23_3_F200_uid1032_bh793_uid1465_In1 <= "" & bh793_w97_11 & bh793_w97_10;
   Compressor_23_3_F200_uid1032_uid1465: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1465_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1465_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1465_Out0_copy1466);
   Compressor_23_3_F200_uid1032_bh793_uid1465_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1465_Out0_copy1466; -- output copy to hold a pipeline register if needed

   bh793_w96_13 <= Compressor_23_3_F200_uid1032_bh793_uid1465_Out0(0);
   bh793_w97_12 <= Compressor_23_3_F200_uid1032_bh793_uid1465_Out0(1);
   bh793_w98_11 <= Compressor_23_3_F200_uid1032_bh793_uid1465_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1467_In0 <= "" & bh793_w98_9 & bh793_w98_10 & "0";
   Compressor_3_2_F200_uid1040_uid1467: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1467_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1467_Out0_copy1468);
   Compressor_3_2_F200_uid1040_bh793_uid1467_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1467_Out0_copy1468; -- output copy to hold a pipeline register if needed

   bh793_w98_12 <= Compressor_3_2_F200_uid1040_bh793_uid1467_Out0(0);
   bh793_w99_12 <= Compressor_3_2_F200_uid1040_bh793_uid1467_Out0(1);

   Compressor_23_3_F200_uid1032_bh793_uid1469_In0 <= "" & bh793_w99_9 & bh793_w99_11 & bh793_w99_10;
   Compressor_23_3_F200_uid1032_bh793_uid1469_In1 <= "" & bh793_w100_9 & bh793_w100_6;
   Compressor_23_3_F200_uid1032_uid1469: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1469_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1469_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1469_Out0_copy1470);
   Compressor_23_3_F200_uid1032_bh793_uid1469_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1469_Out0_copy1470; -- output copy to hold a pipeline register if needed

   bh793_w99_13 <= Compressor_23_3_F200_uid1032_bh793_uid1469_Out0(0);
   bh793_w100_10 <= Compressor_23_3_F200_uid1032_bh793_uid1469_Out0(1);
   bh793_w101_8 <= Compressor_23_3_F200_uid1032_bh793_uid1469_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1471_In0 <= "" & bh793_w101_7 & bh793_w101_6 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1471_In1 <= "" & bh793_w102_7 & bh793_w102_4;
   Compressor_23_3_F200_uid1032_uid1471: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1471_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1471_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1471_Out0_copy1472);
   Compressor_23_3_F200_uid1032_bh793_uid1471_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1471_Out0_copy1472; -- output copy to hold a pipeline register if needed

   bh793_w101_9 <= Compressor_23_3_F200_uid1032_bh793_uid1471_Out0(0);
   bh793_w102_8 <= Compressor_23_3_F200_uid1032_bh793_uid1471_Out0(1);
   bh793_w103_5 <= Compressor_23_3_F200_uid1032_bh793_uid1471_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1473_In0 <= "" & bh793_w103_4 & bh793_w103_3 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1473_In1 <= "" & bh793_w104_2;
   Compressor_14_3_F200_uid1054_uid1473: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1473_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1473_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1473_Out0_copy1474);
   Compressor_14_3_F200_uid1054_bh793_uid1473_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1473_Out0_copy1474; -- output copy to hold a pipeline register if needed

   bh793_w103_6 <= Compressor_14_3_F200_uid1054_bh793_uid1473_Out0(0);
   bh793_w104_3 <= Compressor_14_3_F200_uid1054_bh793_uid1473_Out0(1);
   bh793_w105_2 <= Compressor_14_3_F200_uid1054_bh793_uid1473_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1475_In0 <= "" & bh793_w105_1 & bh793_w105_0 & "0";
   Compressor_3_2_F200_uid1040_uid1475: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1475_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1475_Out0_copy1476);
   Compressor_3_2_F200_uid1040_bh793_uid1475_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1475_Out0_copy1476; -- output copy to hold a pipeline register if needed

   bh793_w105_3 <= Compressor_3_2_F200_uid1040_bh793_uid1475_Out0(0);

   Compressor_14_3_F200_uid1054_bh793_uid1477_In0 <= "" & bh793_w23_7 & bh793_w23_6 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1477_In1 <= "" & bh793_w24_6;
   Compressor_14_3_F200_uid1054_uid1477: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1477_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1477_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1477_Out0_copy1478);
   Compressor_14_3_F200_uid1054_bh793_uid1477_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1477_Out0_copy1478; -- output copy to hold a pipeline register if needed

   bh793_w23_8 <= Compressor_14_3_F200_uid1054_bh793_uid1477_Out0(0);
   bh793_w24_7 <= Compressor_14_3_F200_uid1054_bh793_uid1477_Out0(1);
   bh793_w25_8 <= Compressor_14_3_F200_uid1054_bh793_uid1477_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1479_In0 <= "" & bh793_w25_7 & bh793_w25_6 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1479_In1 <= "" & bh793_w26_6;
   Compressor_14_3_F200_uid1054_uid1479: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1479_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1479_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1479_Out0_copy1480);
   Compressor_14_3_F200_uid1054_bh793_uid1479_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1479_Out0_copy1480; -- output copy to hold a pipeline register if needed

   bh793_w25_9 <= Compressor_14_3_F200_uid1054_bh793_uid1479_Out0(0);
   bh793_w26_7 <= Compressor_14_3_F200_uid1054_bh793_uid1479_Out0(1);
   bh793_w27_8 <= Compressor_14_3_F200_uid1054_bh793_uid1479_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1481_In0 <= "" & bh793_w27_7 & bh793_w27_6 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1481_In1 <= "" & bh793_w28_6;
   Compressor_14_3_F200_uid1054_uid1481: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1481_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1481_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1481_Out0_copy1482);
   Compressor_14_3_F200_uid1054_bh793_uid1481_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1481_Out0_copy1482; -- output copy to hold a pipeline register if needed

   bh793_w27_9 <= Compressor_14_3_F200_uid1054_bh793_uid1481_Out0(0);
   bh793_w28_7 <= Compressor_14_3_F200_uid1054_bh793_uid1481_Out0(1);
   bh793_w29_8 <= Compressor_14_3_F200_uid1054_bh793_uid1481_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1483_In0 <= "" & bh793_w29_7 & bh793_w29_6 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1483_In1 <= "" & bh793_w30_6;
   Compressor_14_3_F200_uid1054_uid1483: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1483_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1483_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1483_Out0_copy1484);
   Compressor_14_3_F200_uid1054_bh793_uid1483_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1483_Out0_copy1484; -- output copy to hold a pipeline register if needed

   bh793_w29_9 <= Compressor_14_3_F200_uid1054_bh793_uid1483_Out0(0);
   bh793_w30_7 <= Compressor_14_3_F200_uid1054_bh793_uid1483_Out0(1);
   bh793_w31_8 <= Compressor_14_3_F200_uid1054_bh793_uid1483_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1485_In0 <= "" & bh793_w31_7 & bh793_w31_6 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1485_In1 <= "" & bh793_w32_6;
   Compressor_14_3_F200_uid1054_uid1485: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1485_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1485_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1485_Out0_copy1486);
   Compressor_14_3_F200_uid1054_bh793_uid1485_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1485_Out0_copy1486; -- output copy to hold a pipeline register if needed

   bh793_w31_9 <= Compressor_14_3_F200_uid1054_bh793_uid1485_Out0(0);
   bh793_w32_7 <= Compressor_14_3_F200_uid1054_bh793_uid1485_Out0(1);
   bh793_w33_8 <= Compressor_14_3_F200_uid1054_bh793_uid1485_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1487_In0 <= "" & bh793_w33_7 & bh793_w33_6 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1487_In1 <= "" & bh793_w34_7;
   Compressor_14_3_F200_uid1054_uid1487: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1487_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1487_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1487_Out0_copy1488);
   Compressor_14_3_F200_uid1054_bh793_uid1487_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1487_Out0_copy1488; -- output copy to hold a pipeline register if needed

   bh793_w33_9 <= Compressor_14_3_F200_uid1054_bh793_uid1487_Out0(0);
   bh793_w34_8 <= Compressor_14_3_F200_uid1054_bh793_uid1487_Out0(1);
   bh793_w35_10 <= Compressor_14_3_F200_uid1054_bh793_uid1487_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1489_In0 <= "" & bh793_w35_9 & bh793_w35_8 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1489_In1 <= "" & bh793_w36_9;
   Compressor_14_3_F200_uid1054_uid1489: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1489_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1489_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1489_Out0_copy1490);
   Compressor_14_3_F200_uid1054_bh793_uid1489_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1489_Out0_copy1490; -- output copy to hold a pipeline register if needed

   bh793_w35_11 <= Compressor_14_3_F200_uid1054_bh793_uid1489_Out0(0);
   bh793_w36_10 <= Compressor_14_3_F200_uid1054_bh793_uid1489_Out0(1);
   bh793_w37_8 <= Compressor_14_3_F200_uid1054_bh793_uid1489_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1491_In0 <= "" & bh793_w37_7 & bh793_w37_6 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1491_In1 <= "" & bh793_w38_9;
   Compressor_14_3_F200_uid1054_uid1491: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1491_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1491_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1491_Out0_copy1492);
   Compressor_14_3_F200_uid1054_bh793_uid1491_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1491_Out0_copy1492; -- output copy to hold a pipeline register if needed

   bh793_w37_9 <= Compressor_14_3_F200_uid1054_bh793_uid1491_Out0(0);
   bh793_w38_10 <= Compressor_14_3_F200_uid1054_bh793_uid1491_Out0(1);
   bh793_w39_8 <= Compressor_14_3_F200_uid1054_bh793_uid1491_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1493_In0 <= "" & bh793_w40_10 & bh793_w40_9 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1493_In1 <= "" & bh793_w41_7;
   Compressor_14_3_F200_uid1054_uid1493: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1493_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1493_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1493_Out0_copy1494);
   Compressor_14_3_F200_uid1054_bh793_uid1493_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1493_Out0_copy1494; -- output copy to hold a pipeline register if needed

   bh793_w40_11 <= Compressor_14_3_F200_uid1054_bh793_uid1493_Out0(0);
   bh793_w41_8 <= Compressor_14_3_F200_uid1054_bh793_uid1493_Out0(1);
   bh793_w42_11 <= Compressor_14_3_F200_uid1054_bh793_uid1493_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1495_In0 <= "" & bh793_w42_10 & bh793_w42_9 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1495_In1 <= "" & bh793_w43_7;
   Compressor_14_3_F200_uid1054_uid1495: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1495_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1495_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1495_Out0_copy1496);
   Compressor_14_3_F200_uid1054_bh793_uid1495_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1495_Out0_copy1496; -- output copy to hold a pipeline register if needed

   bh793_w42_12 <= Compressor_14_3_F200_uid1054_bh793_uid1495_Out0(0);
   bh793_w43_8 <= Compressor_14_3_F200_uid1054_bh793_uid1495_Out0(1);
   bh793_w44_11 <= Compressor_14_3_F200_uid1054_bh793_uid1495_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1497_In0 <= "" & bh793_w44_10 & bh793_w44_9 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1497_In1 <= "" & bh793_w45_7;
   Compressor_14_3_F200_uid1054_uid1497: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1497_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1497_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1497_Out0_copy1498);
   Compressor_14_3_F200_uid1054_bh793_uid1497_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1497_Out0_copy1498; -- output copy to hold a pipeline register if needed

   bh793_w44_12 <= Compressor_14_3_F200_uid1054_bh793_uid1497_Out0(0);
   bh793_w45_8 <= Compressor_14_3_F200_uid1054_bh793_uid1497_Out0(1);
   bh793_w46_11 <= Compressor_14_3_F200_uid1054_bh793_uid1497_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1499_In0 <= "" & bh793_w46_10 & bh793_w46_9 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1499_In1 <= "" & bh793_w47_7;
   Compressor_14_3_F200_uid1054_uid1499: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1499_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1499_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1499_Out0_copy1500);
   Compressor_14_3_F200_uid1054_bh793_uid1499_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1499_Out0_copy1500; -- output copy to hold a pipeline register if needed

   bh793_w46_12 <= Compressor_14_3_F200_uid1054_bh793_uid1499_Out0(0);
   bh793_w47_8 <= Compressor_14_3_F200_uid1054_bh793_uid1499_Out0(1);
   bh793_w48_12 <= Compressor_14_3_F200_uid1054_bh793_uid1499_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1501_In0 <= "" & bh793_w48_11 & bh793_w48_10 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1501_In1 <= "" & bh793_w49_9;
   Compressor_14_3_F200_uid1054_uid1501: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1501_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1501_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1501_Out0_copy1502);
   Compressor_14_3_F200_uid1054_bh793_uid1501_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1501_Out0_copy1502; -- output copy to hold a pipeline register if needed

   bh793_w48_13 <= Compressor_14_3_F200_uid1054_bh793_uid1501_Out0(0);
   bh793_w49_10 <= Compressor_14_3_F200_uid1054_bh793_uid1501_Out0(1);
   bh793_w50_14 <= Compressor_14_3_F200_uid1054_bh793_uid1501_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1503_In0 <= "" & bh793_w50_12 & bh793_w50_13 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1503_In1 <= "" & bh793_w51_12;
   Compressor_14_3_F200_uid1054_uid1503: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1503_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1503_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1503_Out0_copy1504);
   Compressor_14_3_F200_uid1054_bh793_uid1503_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1503_Out0_copy1504; -- output copy to hold a pipeline register if needed

   bh793_w50_15 <= Compressor_14_3_F200_uid1054_bh793_uid1503_Out0(0);
   bh793_w51_13 <= Compressor_14_3_F200_uid1054_bh793_uid1503_Out0(1);
   bh793_w52_18 <= Compressor_14_3_F200_uid1054_bh793_uid1503_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1505_In0 <= "" & bh793_w52_16 & bh793_w52_17 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1505_In1 <= "" & bh793_w53_15;
   Compressor_14_3_F200_uid1054_uid1505: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1505_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1505_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1505_Out0_copy1506);
   Compressor_14_3_F200_uid1054_bh793_uid1505_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1505_Out0_copy1506; -- output copy to hold a pipeline register if needed

   bh793_w52_19 <= Compressor_14_3_F200_uid1054_bh793_uid1505_Out0(0);
   bh793_w53_16 <= Compressor_14_3_F200_uid1054_bh793_uid1505_Out0(1);
   bh793_w54_20 <= Compressor_14_3_F200_uid1054_bh793_uid1505_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1507_In0 <= "" & bh793_w54_18 & bh793_w54_19 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1507_In1 <= "" & bh793_w55_17 & bh793_w55_18;
   Compressor_23_3_F200_uid1032_uid1507: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1507_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1507_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1507_Out0_copy1508);
   Compressor_23_3_F200_uid1032_bh793_uid1507_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1507_Out0_copy1508; -- output copy to hold a pipeline register if needed

   bh793_w54_21 <= Compressor_23_3_F200_uid1032_bh793_uid1507_Out0(0);
   bh793_w55_19 <= Compressor_23_3_F200_uid1032_bh793_uid1507_Out0(1);
   bh793_w56_20 <= Compressor_23_3_F200_uid1032_bh793_uid1507_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1509_In0 <= "" & bh793_w56_18 & bh793_w56_19 & "0";
   Compressor_3_2_F200_uid1040_uid1509: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1509_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1509_Out0_copy1510);
   Compressor_3_2_F200_uid1040_bh793_uid1509_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1509_Out0_copy1510; -- output copy to hold a pipeline register if needed

   bh793_w56_21 <= Compressor_3_2_F200_uid1040_bh793_uid1509_Out0(0);
   bh793_w57_20 <= Compressor_3_2_F200_uid1040_bh793_uid1509_Out0(1);

   Compressor_23_3_F200_uid1032_bh793_uid1511_In0 <= "" & bh793_w57_17 & bh793_w57_18 & bh793_w57_19;
   Compressor_23_3_F200_uid1032_bh793_uid1511_In1 <= "" & bh793_w58_17 & bh793_w58_18;
   Compressor_23_3_F200_uid1032_uid1511: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1511_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1511_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1511_Out0_copy1512);
   Compressor_23_3_F200_uid1032_bh793_uid1511_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1511_Out0_copy1512; -- output copy to hold a pipeline register if needed

   bh793_w57_21 <= Compressor_23_3_F200_uid1032_bh793_uid1511_Out0(0);
   bh793_w58_19 <= Compressor_23_3_F200_uid1032_bh793_uid1511_Out0(1);
   bh793_w59_20 <= Compressor_23_3_F200_uid1032_bh793_uid1511_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1513_In0 <= "" & bh793_w59_18 & bh793_w59_19 & "0";
   Compressor_3_2_F200_uid1040_uid1513: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1513_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1513_Out0_copy1514);
   Compressor_3_2_F200_uid1040_bh793_uid1513_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1513_Out0_copy1514; -- output copy to hold a pipeline register if needed

   bh793_w59_21 <= Compressor_3_2_F200_uid1040_bh793_uid1513_Out0(0);
   bh793_w60_20 <= Compressor_3_2_F200_uid1040_bh793_uid1513_Out0(1);

   Compressor_23_3_F200_uid1032_bh793_uid1515_In0 <= "" & bh793_w60_17 & bh793_w60_18 & bh793_w60_19;
   Compressor_23_3_F200_uid1032_bh793_uid1515_In1 <= "" & bh793_w61_17 & bh793_w61_18;
   Compressor_23_3_F200_uid1032_uid1515: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1515_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1515_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1515_Out0_copy1516);
   Compressor_23_3_F200_uid1032_bh793_uid1515_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1515_Out0_copy1516; -- output copy to hold a pipeline register if needed

   bh793_w60_21 <= Compressor_23_3_F200_uid1032_bh793_uid1515_Out0(0);
   bh793_w61_19 <= Compressor_23_3_F200_uid1032_bh793_uid1515_Out0(1);
   bh793_w62_20 <= Compressor_23_3_F200_uid1032_bh793_uid1515_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1517_In0 <= "" & bh793_w62_18 & bh793_w62_19 & "0";
   Compressor_3_2_F200_uid1040_uid1517: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1517_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1517_Out0_copy1518);
   Compressor_3_2_F200_uid1040_bh793_uid1517_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1517_Out0_copy1518; -- output copy to hold a pipeline register if needed

   bh793_w62_21 <= Compressor_3_2_F200_uid1040_bh793_uid1517_Out0(0);
   bh793_w63_20 <= Compressor_3_2_F200_uid1040_bh793_uid1517_Out0(1);

   Compressor_23_3_F200_uid1032_bh793_uid1519_In0 <= "" & bh793_w63_17 & bh793_w63_18 & bh793_w63_19;
   Compressor_23_3_F200_uid1032_bh793_uid1519_In1 <= "" & bh793_w64_17 & bh793_w64_18;
   Compressor_23_3_F200_uid1032_uid1519: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1519_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1519_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1519_Out0_copy1520);
   Compressor_23_3_F200_uid1032_bh793_uid1519_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1519_Out0_copy1520; -- output copy to hold a pipeline register if needed

   bh793_w63_21 <= Compressor_23_3_F200_uid1032_bh793_uid1519_Out0(0);
   bh793_w64_19 <= Compressor_23_3_F200_uid1032_bh793_uid1519_Out0(1);
   bh793_w65_20 <= Compressor_23_3_F200_uid1032_bh793_uid1519_Out0(2);

   Compressor_3_2_F200_uid1040_bh793_uid1521_In0 <= "" & bh793_w65_18 & bh793_w65_19 & "0";
   Compressor_3_2_F200_uid1040_uid1521: Compressor_3_2_F200_uid1040
      port map ( X0 => Compressor_3_2_F200_uid1040_bh793_uid1521_In0,
                 R => Compressor_3_2_F200_uid1040_bh793_uid1521_Out0_copy1522);
   Compressor_3_2_F200_uid1040_bh793_uid1521_Out0 <= Compressor_3_2_F200_uid1040_bh793_uid1521_Out0_copy1522; -- output copy to hold a pipeline register if needed

   bh793_w65_21 <= Compressor_3_2_F200_uid1040_bh793_uid1521_Out0(0);
   bh793_w66_19 <= Compressor_3_2_F200_uid1040_bh793_uid1521_Out0(1);

   Compressor_23_3_F200_uid1032_bh793_uid1523_In0 <= "" & bh793_w66_16 & bh793_w66_17 & bh793_w66_18;
   Compressor_23_3_F200_uid1032_bh793_uid1523_In1 <= "" & bh793_w67_16 & bh793_w67_15;
   Compressor_23_3_F200_uid1032_uid1523: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1523_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1523_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1523_Out0_copy1524);
   Compressor_23_3_F200_uid1032_bh793_uid1523_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1523_Out0_copy1524; -- output copy to hold a pipeline register if needed

   bh793_w66_20 <= Compressor_23_3_F200_uid1032_bh793_uid1523_Out0(0);
   bh793_w67_17 <= Compressor_23_3_F200_uid1032_bh793_uid1523_Out0(1);
   bh793_w68_19 <= Compressor_23_3_F200_uid1032_bh793_uid1523_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1525_In0 <= "" & bh793_w68_17 & bh793_w68_18 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1525_In1 <= "" & bh793_w69_15 & bh793_w69_12;
   Compressor_23_3_F200_uid1032_uid1525: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1525_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1525_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1525_Out0_copy1526);
   Compressor_23_3_F200_uid1032_bh793_uid1525_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1525_Out0_copy1526; -- output copy to hold a pipeline register if needed

   bh793_w68_20 <= Compressor_23_3_F200_uid1032_bh793_uid1525_Out0(0);
   bh793_w69_16 <= Compressor_23_3_F200_uid1032_bh793_uid1525_Out0(1);
   bh793_w70_18 <= Compressor_23_3_F200_uid1032_bh793_uid1525_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1527_In0 <= "" & bh793_w70_16 & bh793_w70_17 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1527_In1 <= "" & bh793_w71_16 & bh793_w71_14;
   Compressor_23_3_F200_uid1032_uid1527: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1527_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1527_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1527_Out0_copy1528);
   Compressor_23_3_F200_uid1032_bh793_uid1527_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1527_Out0_copy1528; -- output copy to hold a pipeline register if needed

   bh793_w70_19 <= Compressor_23_3_F200_uid1032_bh793_uid1527_Out0(0);
   bh793_w71_17 <= Compressor_23_3_F200_uid1032_bh793_uid1527_Out0(1);
   bh793_w72_17 <= Compressor_23_3_F200_uid1032_bh793_uid1527_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1529_In0 <= "" & bh793_w72_16 & bh793_w72_15 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1529_In1 <= "" & bh793_w73_17 & bh793_w73_16;
   Compressor_23_3_F200_uid1032_uid1529: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1529_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1529_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1529_Out0_copy1530);
   Compressor_23_3_F200_uid1032_bh793_uid1529_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1529_Out0_copy1530; -- output copy to hold a pipeline register if needed

   bh793_w72_18 <= Compressor_23_3_F200_uid1032_bh793_uid1529_Out0(0);
   bh793_w73_18 <= Compressor_23_3_F200_uid1032_bh793_uid1529_Out0(1);
   bh793_w74_17 <= Compressor_23_3_F200_uid1032_bh793_uid1529_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1531_In0 <= "" & bh793_w74_16 & bh793_w74_14 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1531_In1 <= "" & bh793_w75_16 & bh793_w75_15;
   Compressor_23_3_F200_uid1032_uid1531: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1531_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1531_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1531_Out0_copy1532);
   Compressor_23_3_F200_uid1032_bh793_uid1531_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1531_Out0_copy1532; -- output copy to hold a pipeline register if needed

   bh793_w74_18 <= Compressor_23_3_F200_uid1032_bh793_uid1531_Out0(0);
   bh793_w75_17 <= Compressor_23_3_F200_uid1032_bh793_uid1531_Out0(1);
   bh793_w76_18 <= Compressor_23_3_F200_uid1032_bh793_uid1531_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1533_In0 <= "" & bh793_w76_17 & bh793_w76_16 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1533_In1 <= "" & bh793_w77_14 & bh793_w77_12;
   Compressor_23_3_F200_uid1032_uid1533: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1533_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1533_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1533_Out0_copy1534);
   Compressor_23_3_F200_uid1032_bh793_uid1533_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1533_Out0_copy1534; -- output copy to hold a pipeline register if needed

   bh793_w76_19 <= Compressor_23_3_F200_uid1032_bh793_uid1533_Out0(0);
   bh793_w77_15 <= Compressor_23_3_F200_uid1032_bh793_uid1533_Out0(1);
   bh793_w78_16 <= Compressor_23_3_F200_uid1032_bh793_uid1533_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1535_In0 <= "" & bh793_w78_15 & bh793_w78_14 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1535_In1 <= "" & bh793_w79_12 & bh793_w79_10;
   Compressor_23_3_F200_uid1032_uid1535: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1535_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1535_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1535_Out0_copy1536);
   Compressor_23_3_F200_uid1032_bh793_uid1535_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1535_Out0_copy1536; -- output copy to hold a pipeline register if needed

   bh793_w78_17 <= Compressor_23_3_F200_uid1032_bh793_uid1535_Out0(0);
   bh793_w79_13 <= Compressor_23_3_F200_uid1032_bh793_uid1535_Out0(1);
   bh793_w80_17 <= Compressor_23_3_F200_uid1032_bh793_uid1535_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1537_In0 <= "" & bh793_w80_16 & bh793_w80_15 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1537_In1 <= "" & bh793_w81_13;
   Compressor_14_3_F200_uid1054_uid1537: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1537_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1537_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1537_Out0_copy1538);
   Compressor_14_3_F200_uid1054_bh793_uid1537_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1537_Out0_copy1538; -- output copy to hold a pipeline register if needed

   bh793_w80_18 <= Compressor_14_3_F200_uid1054_bh793_uid1537_Out0(0);
   bh793_w81_14 <= Compressor_14_3_F200_uid1054_bh793_uid1537_Out0(1);
   bh793_w82_16 <= Compressor_14_3_F200_uid1054_bh793_uid1537_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1539_In0 <= "" & bh793_w82_15 & bh793_w82_14 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1539_In1 <= "" & bh793_w83_12 & bh793_w83_10;
   Compressor_23_3_F200_uid1032_uid1539: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1539_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1539_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1539_Out0_copy1540);
   Compressor_23_3_F200_uid1032_bh793_uid1539_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1539_Out0_copy1540; -- output copy to hold a pipeline register if needed

   bh793_w82_17 <= Compressor_23_3_F200_uid1032_bh793_uid1539_Out0(0);
   bh793_w83_13 <= Compressor_23_3_F200_uid1032_bh793_uid1539_Out0(1);
   bh793_w84_13 <= Compressor_23_3_F200_uid1032_bh793_uid1539_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1541_In0 <= "" & bh793_w84_12 & bh793_w84_11 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1541_In1 <= "" & bh793_w85_12;
   Compressor_14_3_F200_uid1054_uid1541: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1541_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1541_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1541_Out0_copy1542);
   Compressor_14_3_F200_uid1054_bh793_uid1541_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1541_Out0_copy1542; -- output copy to hold a pipeline register if needed

   bh793_w84_14 <= Compressor_14_3_F200_uid1054_bh793_uid1541_Out0(0);
   bh793_w85_13 <= Compressor_14_3_F200_uid1054_bh793_uid1541_Out0(1);
   bh793_w86_13 <= Compressor_14_3_F200_uid1054_bh793_uid1541_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1543_In0 <= "" & bh793_w86_11 & bh793_w86_12 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1543_In1 <= "" & bh793_w87_12 & bh793_w87_13;
   Compressor_23_3_F200_uid1032_uid1543: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1543_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1543_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1543_Out0_copy1544);
   Compressor_23_3_F200_uid1032_bh793_uid1543_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1543_Out0_copy1544; -- output copy to hold a pipeline register if needed

   bh793_w86_14 <= Compressor_23_3_F200_uid1032_bh793_uid1543_Out0(0);
   bh793_w87_14 <= Compressor_23_3_F200_uid1032_bh793_uid1543_Out0(1);
   bh793_w88_13 <= Compressor_23_3_F200_uid1032_bh793_uid1543_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1545_In0 <= "" & bh793_w89_11 & bh793_w89_12 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1545_In1 <= "" & bh793_w90_12 & bh793_w90_13;
   Compressor_23_3_F200_uid1032_uid1545: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1545_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1545_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1545_Out0_copy1546);
   Compressor_23_3_F200_uid1032_bh793_uid1545_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1545_Out0_copy1546; -- output copy to hold a pipeline register if needed

   bh793_w89_13 <= Compressor_23_3_F200_uid1032_bh793_uid1545_Out0(0);
   bh793_w90_14 <= Compressor_23_3_F200_uid1032_bh793_uid1545_Out0(1);
   bh793_w91_13 <= Compressor_23_3_F200_uid1032_bh793_uid1545_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1547_In0 <= "" & bh793_w92_11 & bh793_w92_12 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1547_In1 <= "" & bh793_w93_12 & bh793_w93_13;
   Compressor_23_3_F200_uid1032_uid1547: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1547_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1547_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1547_Out0_copy1548);
   Compressor_23_3_F200_uid1032_bh793_uid1547_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1547_Out0_copy1548; -- output copy to hold a pipeline register if needed

   bh793_w92_13 <= Compressor_23_3_F200_uid1032_bh793_uid1547_Out0(0);
   bh793_w93_14 <= Compressor_23_3_F200_uid1032_bh793_uid1547_Out0(1);
   bh793_w94_13 <= Compressor_23_3_F200_uid1032_bh793_uid1547_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1549_In0 <= "" & bh793_w95_11 & bh793_w95_12 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1549_In1 <= "" & bh793_w96_12 & bh793_w96_13;
   Compressor_23_3_F200_uid1032_uid1549: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1549_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1549_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1549_Out0_copy1550);
   Compressor_23_3_F200_uid1032_bh793_uid1549_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1549_Out0_copy1550; -- output copy to hold a pipeline register if needed

   bh793_w95_13 <= Compressor_23_3_F200_uid1032_bh793_uid1549_Out0(0);
   bh793_w96_14 <= Compressor_23_3_F200_uid1032_bh793_uid1549_Out0(1);
   bh793_w97_13 <= Compressor_23_3_F200_uid1032_bh793_uid1549_Out0(2);

   Compressor_23_3_F200_uid1032_bh793_uid1551_In0 <= "" & bh793_w98_11 & bh793_w98_12 & "0";
   Compressor_23_3_F200_uid1032_bh793_uid1551_In1 <= "" & bh793_w99_12 & bh793_w99_13;
   Compressor_23_3_F200_uid1032_uid1551: Compressor_23_3_F200_uid1032
      port map ( X0 => Compressor_23_3_F200_uid1032_bh793_uid1551_In0,
                 X1 => Compressor_23_3_F200_uid1032_bh793_uid1551_In1,
                 R => Compressor_23_3_F200_uid1032_bh793_uid1551_Out0_copy1552);
   Compressor_23_3_F200_uid1032_bh793_uid1551_Out0 <= Compressor_23_3_F200_uid1032_bh793_uid1551_Out0_copy1552; -- output copy to hold a pipeline register if needed

   bh793_w98_13 <= Compressor_23_3_F200_uid1032_bh793_uid1551_Out0(0);
   bh793_w99_14 <= Compressor_23_3_F200_uid1032_bh793_uid1551_Out0(1);
   bh793_w100_11 <= Compressor_23_3_F200_uid1032_bh793_uid1551_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1553_In0 <= "" & bh793_w101_8 & bh793_w101_9 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1553_In1 <= "" & bh793_w102_8;
   Compressor_14_3_F200_uid1054_uid1553: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1553_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1553_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1553_Out0_copy1554);
   Compressor_14_3_F200_uid1054_bh793_uid1553_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1553_Out0_copy1554; -- output copy to hold a pipeline register if needed

   bh793_w101_10 <= Compressor_14_3_F200_uid1054_bh793_uid1553_Out0(0);
   bh793_w102_9 <= Compressor_14_3_F200_uid1054_bh793_uid1553_Out0(1);
   bh793_w103_7 <= Compressor_14_3_F200_uid1054_bh793_uid1553_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1555_In0 <= "" & bh793_w103_6 & bh793_w103_5 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1555_In1 <= "" & bh793_w104_3;
   Compressor_14_3_F200_uid1054_uid1555: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1555_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1555_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1555_Out0_copy1556);
   Compressor_14_3_F200_uid1054_bh793_uid1555_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1555_Out0_copy1556; -- output copy to hold a pipeline register if needed

   bh793_w103_8 <= Compressor_14_3_F200_uid1054_bh793_uid1555_Out0(0);
   bh793_w104_4 <= Compressor_14_3_F200_uid1054_bh793_uid1555_Out0(1);
   bh793_w105_4 <= Compressor_14_3_F200_uid1054_bh793_uid1555_Out0(2);

   Compressor_14_3_F200_uid1054_bh793_uid1557_In0 <= "" & bh793_w105_3 & bh793_w105_2 & "0" & "0";
   Compressor_14_3_F200_uid1054_bh793_uid1557_In1 <= "" & "0";
   Compressor_14_3_F200_uid1054_uid1557: Compressor_14_3_F200_uid1054
      port map ( X0 => Compressor_14_3_F200_uid1054_bh793_uid1557_In0,
                 X1 => Compressor_14_3_F200_uid1054_bh793_uid1557_In1,
                 R => Compressor_14_3_F200_uid1054_bh793_uid1557_Out0_copy1558);
   Compressor_14_3_F200_uid1054_bh793_uid1557_Out0 <= Compressor_14_3_F200_uid1054_bh793_uid1557_Out0_copy1558; -- output copy to hold a pipeline register if needed

   bh793_w105_5 <= Compressor_14_3_F200_uid1054_bh793_uid1557_Out0(0);
   tmp_bitheapResult_bh793_24 <= bh793_w24_7 & bh793_w23_8 & bh793_w22_4 & bh793_w21_6 & bh793_w20_3 & bh793_w19_4 & bh793_w18_2 & bh793_w17_2 & bh793_w16_0 & bh793_w15_0 & bh793_w14_0 & bh793_w13_0 & bh793_w12_0 & bh793_w11_0 & bh793_w10_0 & bh793_w9_0 & bh793_w8_0 & bh793_w7_0 & bh793_w6_0 & bh793_w5_0 & bh793_w4_0 & bh793_w3_0 & bh793_w2_0 & bh793_w1_0 & bh793_w0_0;

   bitheapFinalAdd_bh793_In0 <= "0" & bh793_w105_5 & bh793_w104_4 & bh793_w103_7 & bh793_w102_9 & bh793_w101_10 & bh793_w100_10 & bh793_w99_14 & bh793_w98_13 & bh793_w97_12 & bh793_w96_14 & bh793_w95_13 & bh793_w94_12 & bh793_w93_14 & bh793_w92_13 & bh793_w91_12 & bh793_w90_14 & bh793_w89_13 & bh793_w88_12 & bh793_w87_14 & bh793_w86_13 & bh793_w85_13 & bh793_w84_14 & bh793_w83_13 & bh793_w82_17 & bh793_w81_14 & bh793_w80_18 & bh793_w79_13 & bh793_w78_17 & bh793_w77_15 & bh793_w76_19 & bh793_w75_17 & bh793_w74_18 & bh793_w73_18 & bh793_w72_17 & bh793_w71_17 & bh793_w70_18 & bh793_w69_16 & bh793_w68_19 & bh793_w67_17 & bh793_w66_19 & bh793_w65_20 & bh793_w64_19 & bh793_w63_20 & bh793_w62_20 & bh793_w61_19 & bh793_w60_20 & bh793_w59_20 & bh793_w58_19 & bh793_w57_20 & bh793_w56_20 & bh793_w55_19 & bh793_w54_20 & bh793_w53_16 & bh793_w52_18 & bh793_w51_13 & bh793_w50_14 & bh793_w49_10 & bh793_w48_13 & bh793_w47_8 & bh793_w46_12 & bh793_w45_8 & bh793_w44_12 & bh793_w43_8 & bh793_w42_12 & bh793_w41_8 & bh793_w40_11 & bh793_w39_8 & bh793_w38_10 & bh793_w37_9 & bh793_w36_10 & bh793_w35_11 & bh793_w34_8 & bh793_w33_9 & bh793_w32_7 & bh793_w31_9 & bh793_w30_7 & bh793_w29_9 & bh793_w28_7 & bh793_w27_9 & bh793_w26_7 & bh793_w25_9;
   bitheapFinalAdd_bh793_In1 <= "0" & bh793_w105_4 & "0" & bh793_w103_8 & "0" & "0" & bh793_w100_11 & "0" & "0" & bh793_w97_13 & "0" & "0" & bh793_w94_13 & "0" & "0" & bh793_w91_13 & "0" & "0" & bh793_w88_13 & "0" & bh793_w86_14 & "0" & bh793_w84_13 & "0" & bh793_w82_16 & "0" & bh793_w80_17 & "0" & bh793_w78_16 & "0" & bh793_w76_18 & "0" & bh793_w74_17 & "0" & bh793_w72_18 & "0" & bh793_w70_19 & "0" & bh793_w68_20 & "0" & bh793_w66_20 & bh793_w65_21 & "0" & bh793_w63_21 & bh793_w62_21 & "0" & bh793_w60_21 & bh793_w59_21 & "0" & bh793_w57_21 & bh793_w56_21 & "0" & bh793_w54_21 & "0" & bh793_w52_19 & "0" & bh793_w50_15 & "0" & bh793_w48_12 & "0" & bh793_w46_11 & "0" & bh793_w44_11 & "0" & bh793_w42_11 & "0" & "0" & bh793_w39_7 & "0" & bh793_w37_8 & "0" & bh793_w35_10 & "0" & bh793_w33_8 & "0" & bh793_w31_8 & "0" & bh793_w29_8 & "0" & bh793_w27_8 & "0" & bh793_w25_8;
   bitheapFinalAdd_bh793_Cin <= '0';

   bitheapFinalAdd_bh793: IntAdder_82_F200_uid1560
      port map ( clk  => clk,
                 Cin => bitheapFinalAdd_bh793_Cin,
                 X => bitheapFinalAdd_bh793_In0,
                 Y => bitheapFinalAdd_bh793_In1,
                 R => bitheapFinalAdd_bh793_Out);
   bitheapResult_bh793 <= bitheapFinalAdd_bh793_Out(80 downto 0) & tmp_bitheapResult_bh793_24;
   R <= bitheapResult_bh793(105 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                  LeftShifter106_by_max_4095_F200_uid1562
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X S padBit
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter106_by_max_4095_F200_uid1562 is
    port (clk : in std_logic;
          X : in  std_logic_vector(105 downto 0);
          S : in  std_logic_vector(11 downto 0);
          padBit : in  std_logic;
          R : out  std_logic_vector(4200 downto 0)   );
end entity;

architecture arch of LeftShifter106_by_max_4095_F200_uid1562 is
signal ps, ps_d1, ps_d2, ps_d3, ps_d4, ps_d5, ps_d6, ps_d7, ps_d8, ps_d9, ps_d10, ps_d11, ps_d12, ps_d13, ps_d14, ps_d15, ps_d16, ps_d17, ps_d18, ps_d19, ps_d20 :  std_logic_vector(11 downto 0);
signal level0 :  std_logic_vector(105 downto 0);
signal level1 :  std_logic_vector(106 downto 0);
signal level2 :  std_logic_vector(108 downto 0);
signal level3, level3_d1 :  std_logic_vector(112 downto 0);
signal level4 :  std_logic_vector(120 downto 0);
signal level5 :  std_logic_vector(136 downto 0);
signal level6 :  std_logic_vector(168 downto 0);
signal level7, level7_d1, level7_d2 :  std_logic_vector(232 downto 0);
signal level8 :  std_logic_vector(360 downto 0);
signal level9, level9_d1, level9_d2, level9_d3 :  std_logic_vector(616 downto 0);
signal level10 :  std_logic_vector(1128 downto 0);
signal level11, level11_d1, level11_d2, level11_d3, level11_d4, level11_d5, level11_d6, level11_d7, level11_d8, level11_d9, level11_d10, level11_d11, level11_d12, level11_d13, level11_d14 :  std_logic_vector(2152 downto 0);
signal level12 :  std_logic_vector(4200 downto 0);
signal padBit_d1, padBit_d2, padBit_d3, padBit_d4, padBit_d5, padBit_d6, padBit_d7, padBit_d8, padBit_d9, padBit_d10, padBit_d11, padBit_d12, padBit_d13, padBit_d14, padBit_d15, padBit_d16, padBit_d17, padBit_d18, padBit_d19, padBit_d20 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            ps_d1 <=  ps;
            ps_d2 <=  ps_d1;
            ps_d3 <=  ps_d2;
            ps_d4 <=  ps_d3;
            ps_d5 <=  ps_d4;
            ps_d6 <=  ps_d5;
            ps_d7 <=  ps_d6;
            ps_d8 <=  ps_d7;
            ps_d9 <=  ps_d8;
            ps_d10 <=  ps_d9;
            ps_d11 <=  ps_d10;
            ps_d12 <=  ps_d11;
            ps_d13 <=  ps_d12;
            ps_d14 <=  ps_d13;
            ps_d15 <=  ps_d14;
            ps_d16 <=  ps_d15;
            ps_d17 <=  ps_d16;
            ps_d18 <=  ps_d17;
            ps_d19 <=  ps_d18;
            ps_d20 <=  ps_d19;
            level3_d1 <=  level3;
            level7_d1 <=  level7;
            level7_d2 <=  level7_d1;
            level9_d1 <=  level9;
            level9_d2 <=  level9_d1;
            level9_d3 <=  level9_d2;
            level11_d1 <=  level11;
            level11_d2 <=  level11_d1;
            level11_d3 <=  level11_d2;
            level11_d4 <=  level11_d3;
            level11_d5 <=  level11_d4;
            level11_d6 <=  level11_d5;
            level11_d7 <=  level11_d6;
            level11_d8 <=  level11_d7;
            level11_d9 <=  level11_d8;
            level11_d10 <=  level11_d9;
            level11_d11 <=  level11_d10;
            level11_d12 <=  level11_d11;
            level11_d13 <=  level11_d12;
            level11_d14 <=  level11_d13;
            padBit_d1 <=  padBit;
            padBit_d2 <=  padBit_d1;
            padBit_d3 <=  padBit_d2;
            padBit_d4 <=  padBit_d3;
            padBit_d5 <=  padBit_d4;
            padBit_d6 <=  padBit_d5;
            padBit_d7 <=  padBit_d6;
            padBit_d8 <=  padBit_d7;
            padBit_d9 <=  padBit_d8;
            padBit_d10 <=  padBit_d9;
            padBit_d11 <=  padBit_d10;
            padBit_d12 <=  padBit_d11;
            padBit_d13 <=  padBit_d12;
            padBit_d14 <=  padBit_d13;
            padBit_d15 <=  padBit_d14;
            padBit_d16 <=  padBit_d15;
            padBit_d17 <=  padBit_d16;
            padBit_d18 <=  padBit_d17;
            padBit_d19 <=  padBit_d18;
            padBit_d20 <=  padBit_d19;
         end if;
      end process;
   ps<= S;
   level0<= X;
   level1<= level0 & (0 downto 0 => '0') when ps(0)= '1' else     (0 downto 0 => padBit) & level0;
   level2<= level1 & (1 downto 0 => '0') when ps(1)= '1' else     (1 downto 0 => padBit) & level1;
   level3<= level2 & (3 downto 0 => '0') when ps(2)= '1' else     (3 downto 0 => padBit) & level2;
   level4<= level3_d1 & (7 downto 0 => '0') when ps_d1(3)= '1' else     (7 downto 0 => padBit_d1) & level3_d1;
   level5<= level4 & (15 downto 0 => '0') when ps_d1(4)= '1' else     (15 downto 0 => padBit_d1) & level4;
   level6<= level5 & (31 downto 0 => '0') when ps_d1(5)= '1' else     (31 downto 0 => padBit_d1) & level5;
   level7<= level6 & (63 downto 0 => '0') when ps_d1(6)= '1' else     (63 downto 0 => padBit_d1) & level6;
   level8<= level7_d2 & (127 downto 0 => '0') when ps_d3(7)= '1' else     (127 downto 0 => padBit_d3) & level7_d2;
   level9<= level8 & (255 downto 0 => '0') when ps_d3(8)= '1' else     (255 downto 0 => padBit_d3) & level8;
   level10<= level9_d3 & (511 downto 0 => '0') when ps_d6(9)= '1' else     (511 downto 0 => padBit_d6) & level9_d3;
   level11<= level10 & (1023 downto 0 => '0') when ps_d6(10)= '1' else     (1023 downto 0 => padBit_d6) & level10;
   level12<= level11_d14 & (2047 downto 0 => '0') when ps_d20(11)= '1' else     (2047 downto 0 => padBit_d20) & level11_d14;
   R <= level12(4200 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                                   s3fdp
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Ledoux Louis - BSC / UPC
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: S3_x S3_y FTZ EOB
-- Output signals: A EOB_Q isNaN

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity s3fdp is
    port (clk, rst : in std_logic;
          S3_x : in  std_logic_vector(65 downto 0);
          S3_y : in  std_logic_vector(65 downto 0);
          FTZ : in  std_logic;
          EOB : in  std_logic;
          A : out  std_logic_vector(99 downto 0);
          EOB_Q : out  std_logic;
          isNaN : out  std_logic   );
end entity;

architecture arch of s3fdp is
   component IntMultiplier_F200_uid791 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(52 downto 0);
             Y : in  std_logic_vector(52 downto 0);
             R : out  std_logic_vector(105 downto 0)   );
   end component;

   component LeftShifter106_by_max_4095_F200_uid1562 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(105 downto 0);
             S : in  std_logic_vector(11 downto 0);
             padBit : in  std_logic;
             R : out  std_logic_vector(4200 downto 0)   );
   end component;

signal sign_X :  std_logic;
signal sign_Y :  std_logic;
signal sign_M, sign_M_d1, sign_M_d2, sign_M_d3, sign_M_d4, sign_M_d5, sign_M_d6, sign_M_d7, sign_M_d8, sign_M_d9, sign_M_d10, sign_M_d11, sign_M_d12, sign_M_d13, sign_M_d14, sign_M_d15, sign_M_d16, sign_M_d17, sign_M_d18, sign_M_d19, sign_M_d20 :  std_logic;
signal isNaN_X :  std_logic;
signal isNaN_Y :  std_logic;
signal isNaN_M, isNaN_M_d1, isNaN_M_d2, isNaN_M_d3, isNaN_M_d4, isNaN_M_d5, isNaN_M_d6, isNaN_M_d7, isNaN_M_d8, isNaN_M_d9, isNaN_M_d10, isNaN_M_d11, isNaN_M_d12, isNaN_M_d13, isNaN_M_d14, isNaN_M_d15, isNaN_M_d16, isNaN_M_d17, isNaN_M_d18, isNaN_M_d19, isNaN_M_d20 :  std_logic;
signal significand_X :  std_logic_vector(52 downto 0);
signal significand_Y :  std_logic_vector(52 downto 0);
signal significand_product :  std_logic_vector(105 downto 0);
signal scale_X_biased :  std_logic_vector(10 downto 0);
signal scale_Y_biased :  std_logic_vector(10 downto 0);
signal scale_product_twice_biased :  std_logic_vector(11 downto 0);
signal significand_product_cpt1 :  std_logic_vector(105 downto 0);
signal shift_value :  std_logic_vector(11 downto 0);
signal shifted_significand :  std_logic_vector(4200 downto 0);
signal too_small, too_small_d1, too_small_d2, too_small_d3, too_small_d4, too_small_d5, too_small_d6, too_small_d7, too_small_d8, too_small_d9, too_small_d10, too_small_d11, too_small_d12, too_small_d13, too_small_d14, too_small_d15, too_small_d16, too_small_d17, too_small_d18, too_small_d19, too_small_d20 :  std_logic;
signal too_big, too_big_d1, too_big_d2, too_big_d3, too_big_d4, too_big_d5, too_big_d6, too_big_d7, too_big_d8, too_big_d9, too_big_d10, too_big_d11, too_big_d12, too_big_d13, too_big_d14, too_big_d15, too_big_d16, too_big_d17, too_big_d18, too_big_d19, too_big_d20 :  std_logic;
signal ext_summand1c :  std_logic_vector(99 downto 0);
signal not_ftz, not_ftz_d1, not_ftz_d2, not_ftz_d3, not_ftz_d4, not_ftz_d5, not_ftz_d6, not_ftz_d7, not_ftz_d8, not_ftz_d9, not_ftz_d10, not_ftz_d11, not_ftz_d12, not_ftz_d13, not_ftz_d14, not_ftz_d15, not_ftz_d16, not_ftz_d17, not_ftz_d18, not_ftz_d19, not_ftz_d20 :  std_logic;
signal EOB_internal, EOB_internal_d1, EOB_internal_d2, EOB_internal_d3, EOB_internal_d4, EOB_internal_d5, EOB_internal_d6, EOB_internal_d7, EOB_internal_d8, EOB_internal_d9, EOB_internal_d10, EOB_internal_d11, EOB_internal_d12, EOB_internal_d13, EOB_internal_d14, EOB_internal_d15, EOB_internal_d16, EOB_internal_d17, EOB_internal_d18, EOB_internal_d19, EOB_internal_d20, EOB_internal_d21 :  std_logic;
signal not_ftz_sync :  std_logic;
signal carry_0_sync :  std_logic;
signal EOB_internal_delayed :  std_logic;
signal isNaN_M_sync :  std_logic;
signal too_big_sync :  std_logic;
signal isNaN_o, isNaN_o_d1 :  std_logic;
signal isNaN_delayed :  std_logic;
signal carry_0 :  std_logic;
signal summand_0 :  std_logic_vector(99 downto 0);
signal summand_and_carry_0 :  std_logic_vector(100 downto 0);
signal acc_0, acc_0_d1 :  std_logic_vector(100 downto 0);
signal acc_0_q :  std_logic_vector(100 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_M_d1 <=  sign_M;
            sign_M_d2 <=  sign_M_d1;
            sign_M_d3 <=  sign_M_d2;
            sign_M_d4 <=  sign_M_d3;
            sign_M_d5 <=  sign_M_d4;
            sign_M_d6 <=  sign_M_d5;
            sign_M_d7 <=  sign_M_d6;
            sign_M_d8 <=  sign_M_d7;
            sign_M_d9 <=  sign_M_d8;
            sign_M_d10 <=  sign_M_d9;
            sign_M_d11 <=  sign_M_d10;
            sign_M_d12 <=  sign_M_d11;
            sign_M_d13 <=  sign_M_d12;
            sign_M_d14 <=  sign_M_d13;
            sign_M_d15 <=  sign_M_d14;
            sign_M_d16 <=  sign_M_d15;
            sign_M_d17 <=  sign_M_d16;
            sign_M_d18 <=  sign_M_d17;
            sign_M_d19 <=  sign_M_d18;
            sign_M_d20 <=  sign_M_d19;
            isNaN_M_d1 <=  isNaN_M;
            isNaN_M_d2 <=  isNaN_M_d1;
            isNaN_M_d3 <=  isNaN_M_d2;
            isNaN_M_d4 <=  isNaN_M_d3;
            isNaN_M_d5 <=  isNaN_M_d4;
            isNaN_M_d6 <=  isNaN_M_d5;
            isNaN_M_d7 <=  isNaN_M_d6;
            isNaN_M_d8 <=  isNaN_M_d7;
            isNaN_M_d9 <=  isNaN_M_d8;
            isNaN_M_d10 <=  isNaN_M_d9;
            isNaN_M_d11 <=  isNaN_M_d10;
            isNaN_M_d12 <=  isNaN_M_d11;
            isNaN_M_d13 <=  isNaN_M_d12;
            isNaN_M_d14 <=  isNaN_M_d13;
            isNaN_M_d15 <=  isNaN_M_d14;
            isNaN_M_d16 <=  isNaN_M_d15;
            isNaN_M_d17 <=  isNaN_M_d16;
            isNaN_M_d18 <=  isNaN_M_d17;
            isNaN_M_d19 <=  isNaN_M_d18;
            isNaN_M_d20 <=  isNaN_M_d19;
            too_small_d1 <=  too_small;
            too_small_d2 <=  too_small_d1;
            too_small_d3 <=  too_small_d2;
            too_small_d4 <=  too_small_d3;
            too_small_d5 <=  too_small_d4;
            too_small_d6 <=  too_small_d5;
            too_small_d7 <=  too_small_d6;
            too_small_d8 <=  too_small_d7;
            too_small_d9 <=  too_small_d8;
            too_small_d10 <=  too_small_d9;
            too_small_d11 <=  too_small_d10;
            too_small_d12 <=  too_small_d11;
            too_small_d13 <=  too_small_d12;
            too_small_d14 <=  too_small_d13;
            too_small_d15 <=  too_small_d14;
            too_small_d16 <=  too_small_d15;
            too_small_d17 <=  too_small_d16;
            too_small_d18 <=  too_small_d17;
            too_small_d19 <=  too_small_d18;
            too_small_d20 <=  too_small_d19;
            too_big_d1 <=  too_big;
            too_big_d2 <=  too_big_d1;
            too_big_d3 <=  too_big_d2;
            too_big_d4 <=  too_big_d3;
            too_big_d5 <=  too_big_d4;
            too_big_d6 <=  too_big_d5;
            too_big_d7 <=  too_big_d6;
            too_big_d8 <=  too_big_d7;
            too_big_d9 <=  too_big_d8;
            too_big_d10 <=  too_big_d9;
            too_big_d11 <=  too_big_d10;
            too_big_d12 <=  too_big_d11;
            too_big_d13 <=  too_big_d12;
            too_big_d14 <=  too_big_d13;
            too_big_d15 <=  too_big_d14;
            too_big_d16 <=  too_big_d15;
            too_big_d17 <=  too_big_d16;
            too_big_d18 <=  too_big_d17;
            too_big_d19 <=  too_big_d18;
            too_big_d20 <=  too_big_d19;
            not_ftz_d1 <=  not_ftz;
            not_ftz_d2 <=  not_ftz_d1;
            not_ftz_d3 <=  not_ftz_d2;
            not_ftz_d4 <=  not_ftz_d3;
            not_ftz_d5 <=  not_ftz_d4;
            not_ftz_d6 <=  not_ftz_d5;
            not_ftz_d7 <=  not_ftz_d6;
            not_ftz_d8 <=  not_ftz_d7;
            not_ftz_d9 <=  not_ftz_d8;
            not_ftz_d10 <=  not_ftz_d9;
            not_ftz_d11 <=  not_ftz_d10;
            not_ftz_d12 <=  not_ftz_d11;
            not_ftz_d13 <=  not_ftz_d12;
            not_ftz_d14 <=  not_ftz_d13;
            not_ftz_d15 <=  not_ftz_d14;
            not_ftz_d16 <=  not_ftz_d15;
            not_ftz_d17 <=  not_ftz_d16;
            not_ftz_d18 <=  not_ftz_d17;
            not_ftz_d19 <=  not_ftz_d18;
            not_ftz_d20 <=  not_ftz_d19;
            EOB_internal_d1 <=  EOB_internal;
            EOB_internal_d2 <=  EOB_internal_d1;
            EOB_internal_d3 <=  EOB_internal_d2;
            EOB_internal_d4 <=  EOB_internal_d3;
            EOB_internal_d5 <=  EOB_internal_d4;
            EOB_internal_d6 <=  EOB_internal_d5;
            EOB_internal_d7 <=  EOB_internal_d6;
            EOB_internal_d8 <=  EOB_internal_d7;
            EOB_internal_d9 <=  EOB_internal_d8;
            EOB_internal_d10 <=  EOB_internal_d9;
            EOB_internal_d11 <=  EOB_internal_d10;
            EOB_internal_d12 <=  EOB_internal_d11;
            EOB_internal_d13 <=  EOB_internal_d12;
            EOB_internal_d14 <=  EOB_internal_d13;
            EOB_internal_d15 <=  EOB_internal_d14;
            EOB_internal_d16 <=  EOB_internal_d15;
            EOB_internal_d17 <=  EOB_internal_d16;
            EOB_internal_d18 <=  EOB_internal_d17;
            EOB_internal_d19 <=  EOB_internal_d18;
            EOB_internal_d20 <=  EOB_internal_d19;
            EOB_internal_d21 <=  EOB_internal_d20;
         end if;
      end process;
   process(clk, rst)
      begin
         if rst = '1' then
            isNaN_o_d1 <=  '0';
            acc_0_d1 <=  (others => '0');
         elsif clk'event and clk = '1' then
            isNaN_o_d1 <=  isNaN_o;
            acc_0_d1 <=  acc_0;
         end if;
      end process;
--------------------------- sign product processing ---------------------------
   sign_X <= S3_x(64);
   sign_Y <= S3_y(64);
   sign_M <= sign_X xor sign_Y;

---------------------------- NaN product processing ----------------------------
   isNaN_X <= S3_x(65);
   isNaN_Y <= S3_y(65);
   isNaN_M <= isNaN_X or isNaN_Y;

---------------------------- significand processing ----------------------------
   significand_X <= S3_x(63 downto 11);
   significand_Y <= S3_y(63 downto 11);
   significand_product_inst: IntMultiplier_F200_uid791
      port map ( clk  => clk,
                 X => significand_X,
                 Y => significand_Y,
                 R => significand_product);

------------------------------- scale processing -------------------------------
   scale_X_biased <= S3_x(10 downto 0);
   scale_Y_biased <= S3_y(10 downto 0);
   scale_product_twice_biased <= ("0" & scale_X_biased) + ("0" & scale_Y_biased);

--------------------------- pre-shift xoring (cpt1) ---------------------------
   significand_product_cpt1 <= significand_product when sign_M='0' else not(significand_product);

------------------------- significand product shifting -------------------------
   shift_value <= (scale_product_twice_biased) - (1995);
   significand_product_shifter_inst: LeftShifter106_by_max_4095_F200_uid1562
      port map ( clk  => clk,
                 S => shift_value,
                 X => significand_product_cpt1,
                 padBit => sign_M,
                 R => shifted_significand);

-------------- detect too low scale for this specific scratchpad --------------
   too_small <= '1' when (shift_value(11)='1') else '0';

-------------- detect too big scale for this specific scratchpad --------------
   too_big <= '1' when (unsigned(shift_value) > 90 and too_small='0') else '0';

--------------- shifted significand part select to form summand ---------------
   ext_summand1c <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" when too_small_d20='1' else shifted_significand(204 downto 105);
----------------------------- Syncing some signals -----------------------------
   not_ftz <= not FTZ;
   EOB_internal <= EOB;
   not_ftz_sync <= not_ftz_d20;
   carry_0_sync <= sign_M_d20;
   EOB_internal_delayed <= EOB_internal_d21;
   isNaN_M_sync <= isNaN_M_d20;
   too_big_sync <= too_big_d20;

------------------------------ Output isNaN latch ------------------------------
   isNaN_o <= (too_big_sync or isNaN_M_sync or isNaN_delayed) when not_ftz_sync='1' else '0';
   isNaN_delayed <= isNaN_o_d1;

---------------------------- Carry Save Accumulator ----------------------------
   -- DQ logic
   acc_0_q <= acc_0_d1;

   -- sequential addition logic
   carry_0 <= carry_0_sync;
   summand_0 <= ext_summand1c(99 downto 0);
   summand_and_carry_0 <= ("0" & summand_0) + carry_0;
   acc_0 <= (("0" & acc_0_q(99 downto 0)) + summand_and_carry_0) when (not_ftz_sync='1') else
            summand_and_carry_0;

-------------------------------- Output Compose --------------------------------
   A <= acc_0_q(99 downto 0);

   EOB_Q <= EOB_internal_delayed;
   isNaN <= isNaN_delayed;
end architecture;

--------------------------------------------------------------------------------
--                                   PE_S3
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Ledoux Louis - BSC / UPC
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: s3_row_i_A s3_col_j_B C_out SOB EOB
-- Output signals: s3_row_im1_A s3_col_jm1_B SOB_Q EOB_Q C_out_Q

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity PE_S3 is
    port (clk, rst : in std_logic;
          s3_row_i_A : in  std_logic_vector(65 downto 0);
          s3_col_j_B : in  std_logic_vector(65 downto 0);
          C_out : in  std_logic_vector(100 downto 0);
          SOB : in  std_logic;
          EOB : in  std_logic;
          s3_row_im1_A : out  std_logic_vector(65 downto 0);
          s3_col_jm1_B : out  std_logic_vector(65 downto 0);
          SOB_Q : out  std_logic;
          EOB_Q : out  std_logic;
          C_out_Q : out  std_logic_vector(100 downto 0)   );
end entity;

architecture arch of PE_S3 is
   component s3fdp is
      port ( clk, rst : in std_logic;
             S3_x : in  std_logic_vector(65 downto 0);
             S3_y : in  std_logic_vector(65 downto 0);
             FTZ : in  std_logic;
             EOB : in  std_logic;
             A : out  std_logic_vector(99 downto 0);
             EOB_Q : out  std_logic;
             isNaN : out  std_logic   );
   end component;

signal s3_row_i_A_q :  std_logic_vector(65 downto 0);
signal s3_col_j_B_q :  std_logic_vector(65 downto 0);
signal sob_delayed :  std_logic;
signal eob_delayed :  std_logic;
signal mux_C_out, mux_C_out_d1, mux_C_out_d2 :  std_logic_vector(100 downto 0);
signal mux_C_out_HSSD :  std_logic_vector(100 downto 0);
signal isNaN_s3fdp :  std_logic;
signal EOB_s3fdp :  std_logic;
signal A_s3fdp :  std_logic_vector(99 downto 0);
signal s3_row_i_A_d1 :  std_logic_vector(65 downto 0);
signal s3_col_j_B_d1 :  std_logic_vector(65 downto 0);
signal SOB_d1 :  std_logic;
signal EOB_d1 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            mux_C_out_d1 <=  mux_C_out;
            mux_C_out_d2 <=  mux_C_out_d1;
            s3_row_i_A_d1 <=  s3_row_i_A;
            s3_col_j_B_d1 <=  s3_col_j_B;
            SOB_d1 <=  SOB;
            EOB_d1 <=  EOB;
         end if;
      end process;
------------------------ Functional delay z-1 of inputs ------------------------
   s3_row_i_A_q <= s3_row_i_A_d1;
   s3_col_j_B_q <= s3_col_j_B_d1;

------------------------- DQ flip flop for SOB and EOB -------------------------
   sob_delayed <= SOB_d1;
   eob_delayed <= EOB_d1;

----------------------------- Half Speed Sink Down -----------------------------
   with EOB_s3fdp  select  mux_C_out <= 
        (isNaN_s3fdp & A_s3fdp) when '1', 
        C_out when others;
   mux_C_out_HSSD <= mux_C_out_d2;

---------------------------- Instantiates the S3FDP ----------------------------
   s3fdp_inst: s3fdp
      port map ( clk => clk,
                 rst  => rst,
                 EOB => EOB,
                 FTZ => SOB,
                 S3_x => s3_row_i_A,
                 S3_y => s3_col_j_B,
                 A => A_s3fdp,
                 EOB_Q => EOB_s3fdp,
                 isNaN => isNaN_s3fdp);

------------------------- Compose the outputs signals -------------------------
   s3_row_im1_A <= s3_row_i_A_q;
   s3_col_jm1_B <= s3_col_j_B_q;
   SOB_Q <= sob_delayed;
   EOB_Q <= eob_delayed;
   C_out_Q <= mux_C_out_HSSD;
end architecture;

--------------------------------------------------------------------------------
--                            SystolicArrayKernel
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Ledoux Louis - BSC / UPC
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: rowsA colsB SOB EOB
-- Output signals: colsC EOB_Q_o

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity SystolicArrayKernel is
    port (clk, rst : in std_logic;
          rowsA : in  std_logic_vector(527 downto 0);
          colsB : in  std_logic_vector(461 downto 0);
          SOB : in  std_logic;
          EOB : in  std_logic;
          colsC : out  std_logic_vector(706 downto 0);
          EOB_Q_o : out  std_logic   );
end entity;

architecture arch of SystolicArrayKernel is
   component PE_S3 is
      port ( clk, rst : in std_logic;
             s3_row_i_A : in  std_logic_vector(65 downto 0);
             s3_col_j_B : in  std_logic_vector(65 downto 0);
             C_out : in  std_logic_vector(100 downto 0);
             SOB : in  std_logic;
             EOB : in  std_logic;
             s3_row_im1_A : out  std_logic_vector(65 downto 0);
             s3_col_jm1_B : out  std_logic_vector(65 downto 0);
             SOB_Q : out  std_logic;
             EOB_Q : out  std_logic;
             C_out_Q : out  std_logic_vector(100 downto 0)   );
   end component;

type T_2D_LAICPT2_np1_m is array(8 downto 0, 6 downto 0) of std_logic_vector(100 downto 0);
type T_2D_n_mp1 is array(7 downto 0, 7 downto 0) of std_logic_vector(65 downto 0);
type T_2D_np1_m is array(8 downto 0, 6 downto 0) of std_logic_vector(65 downto 0);
type T_2D_np1_m_logic is array(8 downto 0, 6 downto 0) of std_logic;
signal systolic_wires_rows_2D : T_2D_n_mp1;
signal systolic_wires_cols_2D : T_2D_np1_m;
signal systolic_sob_2D : T_2D_np1_m_logic;
signal systolic_eob_2D : T_2D_np1_m_logic;
signal systolic_C_out_2D : T_2D_LAICPT2_np1_m;
begin

----------------- Connect bus of B columns to top edges SA PEs -----------------
   cols_in: for JJ in 0 to 6 generate
      systolic_wires_cols_2D(0,JJ) <= colsB(((JJ+1)*66)-1 downto (JJ*66));
   end generate;

------------------ Connect bus of A rows to left edges SA PEs ------------------
   rows_in: for II in 0 to 7 generate
      systolic_wires_rows_2D(II,0) <= rowsA(((II+1)*66)-1 downto (II*66));
   end generate;

-------------- Connect the Start of Block signals of the TOP PEs --------------
   systolic_sob_2D(0,0) <= SOB;
   sob_1st_row: for JJ in 1 to 6 generate
      systolic_sob_2D(0,JJ) <= systolic_sob_2D(1,JJ-1);
   end generate;

--------------- Connect the End of Block signals of the TOP PEs ---------------
   systolic_eob_2D(0,0) <= EOB;
   eob_1st_row: for JJ in 1 to 6 generate
      systolic_eob_2D(0,JJ) <= systolic_eob_2D(1,JJ-1);
   end generate;

----------- Connect with 0s the input C carry out scheme of TOP PEs -----------
   C_out_input_1st_row: for JJ in 0 to 6 generate
      systolic_C_out_2D(0,JJ) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
   end generate;

------------------------- Connect PEs locally together -------------------------
   rows: for II in 0 to 7 generate
      cols: for JJ in 0 to 6 generate
         PE_ij: PE_S3
            port map ( clk => clk,
                       rst => rst,
                       s3_row_i_A => systolic_wires_rows_2D(II,JJ),
                       s3_col_j_B => systolic_wires_cols_2D(II,JJ),
                       SOB => systolic_sob_2D(II,JJ),
                       SOB_Q => systolic_sob_2D(II+1,JJ),
                       EOB => systolic_eob_2D(II,JJ),
                       EOB_Q => systolic_eob_2D(II+1,JJ),
                       C_out => systolic_C_out_2D(II,JJ),
                       C_out_Q => systolic_C_out_2D(II+1,JJ),
                       s3_row_im1_A => systolic_wires_rows_2D(II,JJ+1),
                       s3_col_jm1_B => systolic_wires_cols_2D(II+1,JJ));
      end generate;
   end generate;

------------------ Connect last row output C to output C bus ------------------
   cols_C_out: for JJ in 0 to 6 generate
      colsC(((JJ+1)*101)-1 downto (JJ*101)) <= systolic_C_out_2D(8,JJ);
   end generate;

------ Connect PE(N-1,M-1) EOB_Q to out world for valid data computation ------
   EOB_Q_o <= systolic_eob_2D(8,6);

end architecture;

--------------------------------------------------------------------------------
--                               SystolicArray
--               (SA_orthogonal_8w7h_ieee_11_52_HSSD_F200_uid2)
-- VHDL generated for VirtexUltrascalePlus @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Ledoux Louis - BSC / UPC
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: rowsA colsB SOB EOB
-- Output signals: colsC EOB_Q_o

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity SystolicArray is
    port (clk, rst : in std_logic;
          rowsA : in  std_logic_vector(511 downto 0);
          colsB : in  std_logic_vector(447 downto 0);
          SOB : in  std_logic;
          EOB : in  std_logic;
          colsC : out  std_logic_vector(447 downto 0);
          EOB_Q_o : out  std_logic   );
end entity;

architecture arch of SystolicArray is
   component Arith_to_S3 is
      port ( clk : in std_logic;
             arith_i : in  std_logic_vector(63 downto 0);
             S3_o : out  std_logic_vector(65 downto 0)   );
   end component;

   component l2a is
      port ( clk : in std_logic;
             A : in  std_logic_vector(99 downto 0);
             isNaN : in  std_logic;
             arith_o : out  std_logic_vector(63 downto 0)   );
   end component;

   component SystolicArrayKernel is
      port ( clk, rst : in std_logic;
             rowsA : in  std_logic_vector(527 downto 0);
             colsB : in  std_logic_vector(461 downto 0);
             SOB : in  std_logic;
             EOB : in  std_logic;
             colsC : out  std_logic_vector(706 downto 0);
             EOB_Q_o : out  std_logic   );
   end component;

type array_M_dense is array(6 downto 0) of std_logic_vector(63 downto 0);
type array_M_s3 is array(6 downto 0) of std_logic_vector(65 downto 0);
type array_N_dense is array(7 downto 0) of std_logic_vector(63 downto 0);
type array_N_s3 is array(7 downto 0) of std_logic_vector(65 downto 0);
signal arith_in_row_0 :  std_logic_vector(63 downto 0);
signal arith_in_row_0_q0 :  std_logic_vector(63 downto 0);
signal arith_in_row_1, arith_in_row_1_d1 :  std_logic_vector(63 downto 0);
signal arith_in_row_1_q1 :  std_logic_vector(63 downto 0);
signal arith_in_row_2, arith_in_row_2_d1, arith_in_row_2_d2 :  std_logic_vector(63 downto 0);
signal arith_in_row_2_q2 :  std_logic_vector(63 downto 0);
signal arith_in_row_3, arith_in_row_3_d1, arith_in_row_3_d2, arith_in_row_3_d3 :  std_logic_vector(63 downto 0);
signal arith_in_row_3_q3 :  std_logic_vector(63 downto 0);
signal arith_in_row_4, arith_in_row_4_d1, arith_in_row_4_d2, arith_in_row_4_d3, arith_in_row_4_d4 :  std_logic_vector(63 downto 0);
signal arith_in_row_4_q4 :  std_logic_vector(63 downto 0);
signal arith_in_row_5, arith_in_row_5_d1, arith_in_row_5_d2, arith_in_row_5_d3, arith_in_row_5_d4, arith_in_row_5_d5 :  std_logic_vector(63 downto 0);
signal arith_in_row_5_q5 :  std_logic_vector(63 downto 0);
signal arith_in_row_6, arith_in_row_6_d1, arith_in_row_6_d2, arith_in_row_6_d3, arith_in_row_6_d4, arith_in_row_6_d5, arith_in_row_6_d6 :  std_logic_vector(63 downto 0);
signal arith_in_row_6_q6 :  std_logic_vector(63 downto 0);
signal arith_in_row_7, arith_in_row_7_d1, arith_in_row_7_d2, arith_in_row_7_d3, arith_in_row_7_d4, arith_in_row_7_d5, arith_in_row_7_d6, arith_in_row_7_d7 :  std_logic_vector(63 downto 0);
signal arith_in_row_7_q7 :  std_logic_vector(63 downto 0);
signal arith_in_col_0 :  std_logic_vector(63 downto 0);
signal arith_in_col_0_q0 :  std_logic_vector(63 downto 0);
signal arith_in_col_1, arith_in_col_1_d1 :  std_logic_vector(63 downto 0);
signal arith_in_col_1_q1 :  std_logic_vector(63 downto 0);
signal arith_in_col_2, arith_in_col_2_d1, arith_in_col_2_d2 :  std_logic_vector(63 downto 0);
signal arith_in_col_2_q2 :  std_logic_vector(63 downto 0);
signal arith_in_col_3, arith_in_col_3_d1, arith_in_col_3_d2, arith_in_col_3_d3 :  std_logic_vector(63 downto 0);
signal arith_in_col_3_q3 :  std_logic_vector(63 downto 0);
signal arith_in_col_4, arith_in_col_4_d1, arith_in_col_4_d2, arith_in_col_4_d3, arith_in_col_4_d4 :  std_logic_vector(63 downto 0);
signal arith_in_col_4_q4 :  std_logic_vector(63 downto 0);
signal arith_in_col_5, arith_in_col_5_d1, arith_in_col_5_d2, arith_in_col_5_d3, arith_in_col_5_d4, arith_in_col_5_d5 :  std_logic_vector(63 downto 0);
signal arith_in_col_5_q5 :  std_logic_vector(63 downto 0);
signal arith_in_col_6, arith_in_col_6_d1, arith_in_col_6_d2, arith_in_col_6_d3, arith_in_col_6_d4, arith_in_col_6_d5, arith_in_col_6_d6 :  std_logic_vector(63 downto 0);
signal arith_in_col_6_q6 :  std_logic_vector(63 downto 0);
signal colsC_LAICPT2 :  std_logic_vector(706 downto 0);
signal SOB_select :  std_logic;
signal SOB_q0 :  std_logic;
signal EOB_select :  std_logic;
signal EOB_q0 :  std_logic;
signal LAICPT2_to_arith :  std_logic_vector(447 downto 0);
signal arith_out_col_out_0, arith_out_col_out_0_d1, arith_out_col_out_0_d2, arith_out_col_out_0_d3, arith_out_col_out_0_d4, arith_out_col_out_0_d5, arith_out_col_out_0_d6 :  std_logic_vector(63 downto 0);
signal arith_out_col_out_0_q6 :  std_logic_vector(63 downto 0);
signal arith_out_col_out_1, arith_out_col_out_1_d1, arith_out_col_out_1_d2, arith_out_col_out_1_d3, arith_out_col_out_1_d4, arith_out_col_out_1_d5 :  std_logic_vector(63 downto 0);
signal arith_out_col_out_1_q5 :  std_logic_vector(63 downto 0);
signal arith_out_col_out_2, arith_out_col_out_2_d1, arith_out_col_out_2_d2, arith_out_col_out_2_d3, arith_out_col_out_2_d4 :  std_logic_vector(63 downto 0);
signal arith_out_col_out_2_q4 :  std_logic_vector(63 downto 0);
signal arith_out_col_out_3, arith_out_col_out_3_d1, arith_out_col_out_3_d2, arith_out_col_out_3_d3 :  std_logic_vector(63 downto 0);
signal arith_out_col_out_3_q3 :  std_logic_vector(63 downto 0);
signal arith_out_col_out_4, arith_out_col_out_4_d1, arith_out_col_out_4_d2 :  std_logic_vector(63 downto 0);
signal arith_out_col_out_4_q2 :  std_logic_vector(63 downto 0);
signal arith_out_col_out_5, arith_out_col_out_5_d1 :  std_logic_vector(63 downto 0);
signal arith_out_col_out_5_q1 :  std_logic_vector(63 downto 0);
signal arith_out_col_out_6 :  std_logic_vector(63 downto 0);
signal arith_out_col_out_6_q0 :  std_logic_vector(63 downto 0);
signal rows_i_arith : array_N_dense;
signal rows_i_s3 :  std_logic_vector(527 downto 0);
signal cols_j_arith : array_M_dense;
signal cols_j_s3 :  std_logic_vector(461 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            arith_in_row_1_d1 <=  arith_in_row_1;
            arith_in_row_2_d1 <=  arith_in_row_2;
            arith_in_row_2_d2 <=  arith_in_row_2_d1;
            arith_in_row_3_d1 <=  arith_in_row_3;
            arith_in_row_3_d2 <=  arith_in_row_3_d1;
            arith_in_row_3_d3 <=  arith_in_row_3_d2;
            arith_in_row_4_d1 <=  arith_in_row_4;
            arith_in_row_4_d2 <=  arith_in_row_4_d1;
            arith_in_row_4_d3 <=  arith_in_row_4_d2;
            arith_in_row_4_d4 <=  arith_in_row_4_d3;
            arith_in_row_5_d1 <=  arith_in_row_5;
            arith_in_row_5_d2 <=  arith_in_row_5_d1;
            arith_in_row_5_d3 <=  arith_in_row_5_d2;
            arith_in_row_5_d4 <=  arith_in_row_5_d3;
            arith_in_row_5_d5 <=  arith_in_row_5_d4;
            arith_in_row_6_d1 <=  arith_in_row_6;
            arith_in_row_6_d2 <=  arith_in_row_6_d1;
            arith_in_row_6_d3 <=  arith_in_row_6_d2;
            arith_in_row_6_d4 <=  arith_in_row_6_d3;
            arith_in_row_6_d5 <=  arith_in_row_6_d4;
            arith_in_row_6_d6 <=  arith_in_row_6_d5;
            arith_in_row_7_d1 <=  arith_in_row_7;
            arith_in_row_7_d2 <=  arith_in_row_7_d1;
            arith_in_row_7_d3 <=  arith_in_row_7_d2;
            arith_in_row_7_d4 <=  arith_in_row_7_d3;
            arith_in_row_7_d5 <=  arith_in_row_7_d4;
            arith_in_row_7_d6 <=  arith_in_row_7_d5;
            arith_in_row_7_d7 <=  arith_in_row_7_d6;
            arith_in_col_1_d1 <=  arith_in_col_1;
            arith_in_col_2_d1 <=  arith_in_col_2;
            arith_in_col_2_d2 <=  arith_in_col_2_d1;
            arith_in_col_3_d1 <=  arith_in_col_3;
            arith_in_col_3_d2 <=  arith_in_col_3_d1;
            arith_in_col_3_d3 <=  arith_in_col_3_d2;
            arith_in_col_4_d1 <=  arith_in_col_4;
            arith_in_col_4_d2 <=  arith_in_col_4_d1;
            arith_in_col_4_d3 <=  arith_in_col_4_d2;
            arith_in_col_4_d4 <=  arith_in_col_4_d3;
            arith_in_col_5_d1 <=  arith_in_col_5;
            arith_in_col_5_d2 <=  arith_in_col_5_d1;
            arith_in_col_5_d3 <=  arith_in_col_5_d2;
            arith_in_col_5_d4 <=  arith_in_col_5_d3;
            arith_in_col_5_d5 <=  arith_in_col_5_d4;
            arith_in_col_6_d1 <=  arith_in_col_6;
            arith_in_col_6_d2 <=  arith_in_col_6_d1;
            arith_in_col_6_d3 <=  arith_in_col_6_d2;
            arith_in_col_6_d4 <=  arith_in_col_6_d3;
            arith_in_col_6_d5 <=  arith_in_col_6_d4;
            arith_in_col_6_d6 <=  arith_in_col_6_d5;
            arith_out_col_out_0_d1 <=  arith_out_col_out_0;
            arith_out_col_out_0_d2 <=  arith_out_col_out_0_d1;
            arith_out_col_out_0_d3 <=  arith_out_col_out_0_d2;
            arith_out_col_out_0_d4 <=  arith_out_col_out_0_d3;
            arith_out_col_out_0_d5 <=  arith_out_col_out_0_d4;
            arith_out_col_out_0_d6 <=  arith_out_col_out_0_d5;
            arith_out_col_out_1_d1 <=  arith_out_col_out_1;
            arith_out_col_out_1_d2 <=  arith_out_col_out_1_d1;
            arith_out_col_out_1_d3 <=  arith_out_col_out_1_d2;
            arith_out_col_out_1_d4 <=  arith_out_col_out_1_d3;
            arith_out_col_out_1_d5 <=  arith_out_col_out_1_d4;
            arith_out_col_out_2_d1 <=  arith_out_col_out_2;
            arith_out_col_out_2_d2 <=  arith_out_col_out_2_d1;
            arith_out_col_out_2_d3 <=  arith_out_col_out_2_d2;
            arith_out_col_out_2_d4 <=  arith_out_col_out_2_d3;
            arith_out_col_out_3_d1 <=  arith_out_col_out_3;
            arith_out_col_out_3_d2 <=  arith_out_col_out_3_d1;
            arith_out_col_out_3_d3 <=  arith_out_col_out_3_d2;
            arith_out_col_out_4_d1 <=  arith_out_col_out_4;
            arith_out_col_out_4_d2 <=  arith_out_col_out_4_d1;
            arith_out_col_out_5_d1 <=  arith_out_col_out_5;
         end if;
      end process;
------------ Delay depending on row index incoming dense arithmetic ------------
   arith_in_row_0 <= rowsA(63 downto 0);
   arith_in_row_0_q0 <= arith_in_row_0;
   arith_in_row_1 <= rowsA(127 downto 64);
   arith_in_row_1_q1 <= arith_in_row_1_d1;
   arith_in_row_2 <= rowsA(191 downto 128);
   arith_in_row_2_q2 <= arith_in_row_2_d2;
   arith_in_row_3 <= rowsA(255 downto 192);
   arith_in_row_3_q3 <= arith_in_row_3_d3;
   arith_in_row_4 <= rowsA(319 downto 256);
   arith_in_row_4_q4 <= arith_in_row_4_d4;
   arith_in_row_5 <= rowsA(383 downto 320);
   arith_in_row_5_q5 <= arith_in_row_5_d5;
   arith_in_row_6 <= rowsA(447 downto 384);
   arith_in_row_6_q6 <= arith_in_row_6_d6;
   arith_in_row_7 <= rowsA(511 downto 448);
   arith_in_row_7_q7 <= arith_in_row_7_d7;

------------ Delay depending on col index incoming dense arithmetic ------------
   arith_in_col_0 <= colsB(63 downto 0);
   arith_in_col_0_q0 <= arith_in_col_0;
   arith_in_col_1 <= colsB(127 downto 64);
   arith_in_col_1_q1 <= arith_in_col_1_d1;
   arith_in_col_2 <= colsB(191 downto 128);
   arith_in_col_2_q2 <= arith_in_col_2_d2;
   arith_in_col_3 <= colsB(255 downto 192);
   arith_in_col_3_q3 <= arith_in_col_3_d3;
   arith_in_col_4 <= colsB(319 downto 256);
   arith_in_col_4_q4 <= arith_in_col_4_d4;
   arith_in_col_5 <= colsB(383 downto 320);
   arith_in_col_5_q5 <= arith_in_col_5_d5;
   arith_in_col_6 <= colsB(447 downto 384);
   arith_in_col_6_q6 <= arith_in_col_6_d6;

--------------- Delay SOB/EOB with Arith_to_S3 delay to feed SAK ---------------
   SOB_select <= SOB;
   SOB_q0 <= SOB_select;
   EOB_select <= EOB;
   EOB_q0 <= EOB_select;

--------------- Delay outgoing arithmetic depending on col index ---------------
   arith_out_col_out_0 <= LAICPT2_to_arith(63 downto 0);
   arith_out_col_out_0_q6 <= arith_out_col_out_0_d6;
   arith_out_col_out_1 <= LAICPT2_to_arith(127 downto 64);
   arith_out_col_out_1_q5 <= arith_out_col_out_1_d5;
   arith_out_col_out_2 <= LAICPT2_to_arith(191 downto 128);
   arith_out_col_out_2_q4 <= arith_out_col_out_2_d4;
   arith_out_col_out_3 <= LAICPT2_to_arith(255 downto 192);
   arith_out_col_out_3_q3 <= arith_out_col_out_3_d3;
   arith_out_col_out_4 <= LAICPT2_to_arith(319 downto 256);
   arith_out_col_out_4_q2 <= arith_out_col_out_4_d2;
   arith_out_col_out_5 <= LAICPT2_to_arith(383 downto 320);
   arith_out_col_out_5_q1 <= arith_out_col_out_5_d1;
   arith_out_col_out_6 <= LAICPT2_to_arith(447 downto 384);
   arith_out_col_out_6_q0 <= arith_out_col_out_6;

---------------- Generate Arith_to_S3 for rows and connect them ----------------
   rows_i_arith(0) <= arith_in_row_0_q0;
   rows_i_arith(1) <= arith_in_row_1_q1;
   rows_i_arith(2) <= arith_in_row_2_q2;
   rows_i_arith(3) <= arith_in_row_3_q3;
   rows_i_arith(4) <= arith_in_row_4_q4;
   rows_i_arith(5) <= arith_in_row_5_q5;
   rows_i_arith(6) <= arith_in_row_6_q6;
   rows_i_arith(7) <= arith_in_row_7_q7;
   rows_a2s3: for II in 0 to 7 generate
      a2s3_i: Arith_to_S3
         port map ( clk => clk,
                    arith_i => rows_i_arith(II),
                    s3_o => rows_i_s3(((II+1)*66)-1 downto II*66));
   end generate;

---------------- Generate Arith_to_S3 for cols and connect them ----------------
   cols_j_arith(0) <= arith_in_col_0_q0;
   cols_j_arith(1) <= arith_in_col_1_q1;
   cols_j_arith(2) <= arith_in_col_2_q2;
   cols_j_arith(3) <= arith_in_col_3_q3;
   cols_j_arith(4) <= arith_in_col_4_q4;
   cols_j_arith(5) <= arith_in_col_5_q5;
   cols_j_arith(6) <= arith_in_col_6_q6;
   cols_a2s3: for JJ in 0 to 6 generate
      a2s3_j: Arith_to_S3
         port map ( clk => clk,
                    arith_i => cols_j_arith(JJ),
                    s3_o => cols_j_s3(((JJ+1)*66)-1 downto JJ*66));
   end generate;

-------------------- Instantiate the Systolic Array Kernel --------------------
   sak: SystolicArrayKernel
      port map ( clk => clk,
                 rst => rst,
                 rowsA => rows_i_s3,
                 colsB => cols_j_s3,
                 SOB => SOB_q0,
                 EOB => EOB_q0,
                 EOB_Q_o => EOB_Q_o,
                 colsC => colsC_LAICPT2 );

-------------------------- Generate LAICPT2_to_arith --------------------------
   cols_l2a: for JJ in 0 to 6 generate
      l2a_i: l2a
         port map ( clk => clk,
                    A => colsC_LAICPT2(((JJ+1)*101)-1-1-0 downto JJ*101),
                    isNaN => colsC_LAICPT2(((JJ+1)*101)- 1),
                    arith_o => LAICPT2_to_arith(((JJ+1)*64)-1 downto JJ*64));
   end generate;

-------- Connect outgoing delayed dense arith words to colsC output bus --------
   colsC(63 downto 0) <= arith_out_col_out_0_q6;
   colsC(127 downto 64) <= arith_out_col_out_1_q5;
   colsC(191 downto 128) <= arith_out_col_out_2_q4;
   colsC(255 downto 192) <= arith_out_col_out_3_q3;
   colsC(319 downto 256) <= arith_out_col_out_4_q2;
   colsC(383 downto 320) <= arith_out_col_out_5_q1;
   colsC(447 downto 384) <= arith_out_col_out_6_q0;

end architecture;

